module project2(a,b,opcode,beqout,flow,out);
	wire [31:0] cout;
	wire set,fout;
	input[31:0] a,b;
	input[2:0] opcode;
	output[31:0] out;
	output flow,beqout;
	alu_1 alu0(a[0],b[0],opcode[2],set,opcode,out[0],cout[0]);
	alu_1 alu1(a[1],b[1],cout[0],0,opcode,out[1],cout[1]);
	alu_1 alu2(a[2],b[2],cout[1],0,opcode,out[2],cout[2]);
	alu_1 alu3(a[3],b[3],cout[2],0,opcode,out[3],cout[3]);
	alu_1 alu4(a[4],b[4],cout[3],0,opcode,out[4],cout[4]);
	alu_1 alu5(a[5],b[5],cout[4],0,opcode,out[5],cout[5]);
	alu_1 alu6(a[6],b[6],cout[5],0,opcode,out[6],cout[6]);
	alu_1 alu7(a[7],b[7],cout[6],0,opcode,out[7],cout[7]);
	alu_1 alu8(a[8],b[8],cout[7],0,opcode,out[8],cout[8]);
	alu_1 alu9(a[9],b[9],cout[8],0,opcode,out[9],cout[9]);
	alu_1 alu10(a[10],b[10],cout[9],0,opcode,out[10],cout[10]);
	alu_1 alu11(a[11],b[11],cout[10],0,opcode,out[11],cout[11]);
	alu_1 alu12(a[12],b[12],cout[11],0,opcode,out[12],cout[12]);
	alu_1 alu13(a[13],b[13],cout[12],0,opcode,out[13],cout[13]);
	alu_1 alu14(a[14],b[14],cout[13],0,opcode,out[14],cout[14]);
	alu_1 alu15(a[15],b[15],cout[14],0,opcode,out[15],cout[15]);
	alu_1 alu16(a[16],b[16],cout[15],0,opcode,out[16],cout[16]);
	alu_1 alu17(a[17],b[17],cout[16],0,opcode,out[17],cout[17]);
	alu_1 alu18(a[18],b[18],cout[17],0,opcode,out[18],cout[18]);
	alu_1 alu19(a[19],b[19],cout[18],0,opcode,out[19],cout[19]);
	alu_1 alu20(a[20],b[20],cout[19],0,opcode,out[20],cout[20]);
	alu_1 alu21(a[21],b[21],cout[20],0,opcode,out[21],cout[21]);
	alu_1 alu22(a[22],b[22],cout[21],0,opcode,out[22],cout[22]);
	alu_1 alu23(a[23],b[23],cout[22],0,opcode,out[23],cout[23]);
	alu_1 alu24(a[24],b[24],cout[23],0,opcode,out[24],cout[24]);
	alu_1 alu25(a[25],b[25],cout[24],0,opcode,out[25],cout[25]);
	alu_1 alu26(a[26],b[26],cout[25],0,opcode,out[26],cout[26]);
	alu_1 alu27(a[27],b[27],cout[26],0,opcode,out[27],cout[27]);
	alu_1 alu28(a[28],b[28],cout[27],0,opcode,out[28],cout[28]);
	alu_1 alu29(a[29],b[29],cout[28],0,opcode,out[29],cout[29]);
	alu_1 alu30(a[30],b[30],cout[29],0,opcode,out[30],cout[30]);
	alu_2 alu(a[31],b[31],cout[30],0,opcode,out[31],flow,set);
	or #1
		o(fout,out[0],out[1],out[2],out[3],out[4],out[5],out[6],out[7],out[8],out[9],out[10],out[11],out[12],out[13],out[14],out[15],out[16],out[17],out[18],out[19],out[20],out[21],out[22],out[23],out[24],out[25],out[26],out[27],out[28],out[29],out[30],out[31]);
	not #1
		no(beqout,fout);
	

endmodule
module alu_1(a,b,cin,less,opcode,out,cout);
	input[2:0] opcode;
	input a,b,cin,less;
	output out,cout;
	wire w1,w2,w3,w4,w5;
	wire[2:0] newOP;
	and #1
		a1(w1,a,b);
	or #1
		o1(w2,a,b);
	not #1
		no(w3,b);
	convertBeq convert(newOP,opcode);
	Smallmux submux(w4,newOP[2],b,w3);
	adder add(a,w4,w5,cout,cin);
	Bigmux bm(out,newOP[1:0],w1,w2,w5,less);
		
endmodule
module alu_2(a,b,cin,less,opcode,out,flow,set);
	input[2:0] opcode;
	input a,b,cin,less;
	output out,flow,set;
	wire w1,w2,w3,w4,w5,cout,binvert;
	wire[2:0] newOP;
	and #1
		a1(w1,a,b);
	or #1
		o1(w2,a,b);
	not #1
		no(w3,b);
	convertBeq convert(newOP,opcode);
	Smallmux submux(w4,newOP[2],b,w3);
	adder add(a,w4,w5,cout,cin);
	Bigmux bm(out,newOP[1:0],w1,w2,w5,less);
	xor #1
		xo(flow,cout,cin),
		xo2(set,w5,flow);
endmodule
module adder(a,b,s,cout,cin);
	input a,b,cin;
	output s,cout;
	wire w1,w2,w3,w4; 
	xor #1
		g1(w1,a,b),
		g2(s,w1,cin);
	and #1
		g3(w2,cin,b),
		g4(w3,cin,a),
		g5(w4,a,b);
	or #1
		g6(cout, w2,w3,w4);
endmodule
module Smallmux(cout,opcode,a,b);
	output cout;
	input opcode,a,b;
	wire w1,w2,w3;
	not #1 n1(w1,opcode);
	and #1
		a1(w2,w1,a),
		a2(w3,opcode,b);
	or #1
		o1(cout,w2,w3);
		
endmodule
module Bigmux(cout,opcode,a,b,c,d);
	input[1:0] opcode;
	input a,b,c,d;
	output cout;
	wire w1,w2,w3,w4,w5,w6;
	not #1
		n1(w1,opcode[0]),
		n2(w2,opcode[1]);
	and #1
		a1(w3,w1,w2,a),
		a2(w4,opcode[0],w2,b),
		a3(w5,w1,opcode[1],c),
		a4(w6,opcode[0],opcode[1],d);
	or #1
		o1(cout,w3,w4,w5,w6);
endmodule
module convertBeq(cout,opcode);
	input[2:0] opcode;
	output[2:0] cout;
	or #1 o1(cout[1],opcode[1],opcode[2]);
	and #1
		a1(cout[0],opcode[0],1'b1),
		a2(cout[2],opcode[2],1'b1);
endmodule
	
module test(a,b,opcode,beqout,flow,out); 
	input signed[31:0] out;
	input flow,beqout;
	output [31:0] a,b;
	output[2:0] opcode;
	reg[2:0] opcode;
	reg signed[31:0] a,b;
	project2 alu_32(a,b,opcode,beqout,flow,out);
		
	initial begin
		$monitor($time,,"a=%d b=%d opcode=%b out=%d flow=%d beqout=%d",a,b,opcode,out,flow,beqout);
			#100	a=534924;b=-226972;opcode=100;
			#100	a=-537137;b=3699;opcode=000;
			#100	a=-252140;b=763954;opcode=111;
			#100	a=298145;b=-478283;opcode=000;
			#100	a=-805068;b=303362;opcode=111;
			#100	a=-976767;b=44317;opcode=111;
			#100	a=-234181;b=286003;opcode=100;
			#100	a=418316;b=85201;opcode=111;
			#100	a=714794;b=83346;opcode=010;
			#100	a=232610;b=425822;opcode=100;
			#100	a=-940141;b=-177294;opcode=001;
			#100	a=411026;b=-434494;opcode=001;
			#100	a=-655398;b=312422;opcode=111;
			#100	a=193630;b=-583128;opcode=000;
			#100	a=-965825;b=249368;opcode=010;
			#100	a=-180808;b=119885;opcode=110;
			#100	a=1811;b=-423936;opcode=111;
			#100	a=33020;b=-112010;opcode=001;
			#100	a=331996;b=-288784;opcode=001;
			#100	a=274353;b=794709;opcode=010;
			#100	a=-808062;b=119620;opcode=010;
			#100	a=-535617;b=671005;opcode=110;
			#100	a=-220516;b=937642;opcode=111;
			#100	a=725269;b=-379488;opcode=111;
			#100	a=-930896;b=107901;opcode=001;
			#100	a=-577648;b=906366;opcode=000;
			#100	a=-768343;b=527784;opcode=000;
			#100	a=387514;b=-394783;opcode=100;
			#100	a=-659520;b=-511857;opcode=100;
			#100	a=74155;b=-63636;opcode=000;
			#100	a=223110;b=403067;opcode=111;
			#100	a=-611268;b=-805020;opcode=000;
			#100	a=910183;b=-107126;opcode=000;
			#100	a=279857;b=-263216;opcode=010;
			#100	a=-476842;b=-696091;opcode=111;
			#100	a=-879984;b=498591;opcode=001;
			#100	a=-430831;b=345186;opcode=100;
			#100	a=668842;b=209247;opcode=100;
			#100	a=961329;b=475240;opcode=010;
			#100	a=-358121;b=-217812;opcode=110;
			#100	a=27138;b=-519635;opcode=000;
			#100	a=26025;b=144053;opcode=000;
			#100	a=877886;b=121582;opcode=010;
			#100	a=898020;b=324269;opcode=111;
			#100	a=-175974;b=538622;opcode=001;
			#100	a=308538;b=24295;opcode=111;
			#100	a=738856;b=-937874;opcode=110;
			#100	a=-571508;b=-117128;opcode=111;
			#100	a=-317490;b=-744105;opcode=010;
			#100	a=742209;b=-334022;opcode=111;
			#100	a=-154534;b=129275;opcode=000;
			#100	a=-434032;b=-726519;opcode=001;
			#100	a=-843837;b=-441779;opcode=111;
			#100	a=220377;b=130286;opcode=111;
			#100	a=-247747;b=65022;opcode=111;
			#100	a=-314737;b=-306638;opcode=110;
			#100	a=-728563;b=908054;opcode=000;
			#100	a=209479;b=547457;opcode=100;
			#100	a=-676844;b=-72861;opcode=111;
			#100	a=517879;b=-34233;opcode=110;
			#100	a=-901084;b=565512;opcode=111;
			#100	a=-135650;b=-331057;opcode=110;
			#100	a=-676507;b=-23738;opcode=100;
			#100	a=729023;b=-642184;opcode=110;
			#100	a=707674;b=-906401;opcode=111;
			#100	a=-770711;b=-599339;opcode=100;
			#100	a=-988782;b=-699622;opcode=111;
			#100	a=-756936;b=731360;opcode=110;
			#100	a=-498796;b=465559;opcode=000;
			#100	a=-123313;b=-265600;opcode=010;
			#100	a=-755763;b=705458;opcode=111;
			#100	a=-583383;b=-666937;opcode=110;
			#100	a=529930;b=-461746;opcode=001;
			#100	a=596190;b=341343;opcode=000;
			#100	a=-970821;b=461831;opcode=001;
			#100	a=644410;b=-891242;opcode=001;
			#100	a=633268;b=-15611;opcode=110;
			#100	a=899147;b=-133319;opcode=111;
			#100	a=47119;b=821672;opcode=100;
			#100	a=-204354;b=399433;opcode=100;
			#100	a=-157516;b=157550;opcode=001;
			#100	a=410826;b=-344213;opcode=100;
			#100	a=-788125;b=404862;opcode=111;
			#100	a=-819927;b=-722852;opcode=111;
			#100	a=333748;b=-672892;opcode=110;
			#100	a=155358;b=-330801;opcode=110;
			#100	a=558251;b=159624;opcode=110;
			#100	a=656599;b=327469;opcode=010;
			#100	a=117756;b=709913;opcode=110;
			#100	a=972449;b=-775543;opcode=110;
			#100	a=787762;b=-924855;opcode=010;
			#100	a=652903;b=-683947;opcode=111;
			#100	a=734886;b=948331;opcode=001;
			#100	a=-979400;b=-266950;opcode=100;
			#100	a=-930604;b=-969166;opcode=001;
			#100	a=-416730;b=830362;opcode=100;
			#100	a=435388;b=-633210;opcode=111;
			#100	a=-675506;b=234062;opcode=001;
			#100	a=268323;b=-832170;opcode=001;
			#100	a=-786737;b=-189292;opcode=010;
			#100	a=-882381;b=866238;opcode=110;
			#100	a=879226;b=-625627;opcode=001;
			#100	a=183664;b=743072;opcode=001;
			#100	a=977434;b=146149;opcode=100;
			#100	a=529104;b=210176;opcode=100;
			#100	a=907811;b=-618485;opcode=110;
			#100	a=-966096;b=649822;opcode=111;
			#100	a=670207;b=-60837;opcode=110;
			#100	a=-317732;b=-503601;opcode=000;
			#100	a=-162239;b=930212;opcode=000;
			#100	a=476256;b=843289;opcode=001;
			#100	a=-669685;b=-293239;opcode=100;
			#100	a=-914210;b=887225;opcode=100;
			#100	a=392741;b=866199;opcode=010;
			#100	a=350816;b=-315353;opcode=010;
			#100	a=-576201;b=-415121;opcode=110;
			#100	a=201881;b=-551788;opcode=110;
			#100	a=-140184;b=-235391;opcode=111;
			#100	a=296237;b=200329;opcode=001;
			#100	a=79322;b=-974047;opcode=100;
			#100	a=930187;b=-746223;opcode=010;
			#100	a=-355663;b=-410612;opcode=010;
			#100	a=294219;b=197536;opcode=001;
			#100	a=885174;b=-536480;opcode=010;
			#100	a=314115;b=-527353;opcode=001;
			#100	a=547602;b=-295776;opcode=110;
			#100	a=328962;b=-141784;opcode=111;
			#100	a=899306;b=-666100;opcode=100;
			#100	a=-274020;b=-650964;opcode=001;
			#100	a=-366424;b=-891937;opcode=000;
			#100	a=-197390;b=-835632;opcode=010;
			#100	a=176148;b=-80426;opcode=110;
			#100	a=-205415;b=901197;opcode=010;
			#100	a=24917;b=220255;opcode=000;
			#100	a=-101595;b=897601;opcode=010;
			#100	a=-943227;b=146874;opcode=010;
			#100	a=-320423;b=362394;opcode=111;
			#100	a=258287;b=90818;opcode=110;
			#100	a=-690820;b=833218;opcode=010;
			#100	a=-6313;b=229503;opcode=000;
			#100	a=325573;b=-22491;opcode=110;
			#100	a=206711;b=-502623;opcode=010;
			#100	a=-127001;b=-231025;opcode=111;
			#100	a=-974493;b=-564466;opcode=111;
			#100	a=994016;b=457312;opcode=010;
			#100	a=-35937;b=-566399;opcode=000;
			#100	a=338334;b=51457;opcode=000;
			#100	a=963320;b=328533;opcode=001;
			#100	a=-70885;b=914863;opcode=100;
			#100	a=-100067;b=-416403;opcode=010;
			#100	a=65746;b=417561;opcode=000;
			#100	a=67955;b=-666710;opcode=111;
			#100	a=250820;b=30196;opcode=000;
			#100	a=799459;b=574155;opcode=000;
			#100	a=-309214;b=2020;opcode=110;
			#100	a=555674;b=-562886;opcode=000;
			#100	a=858452;b=-119715;opcode=001;
			#100	a=-632936;b=-438959;opcode=110;
			#100	a=800871;b=-936407;opcode=111;
			#100	a=-924824;b=166450;opcode=111;
			#100	a=-502029;b=283522;opcode=110;
			#100	a=635052;b=905617;opcode=000;
			#100	a=732289;b=-842367;opcode=000;
			#100	a=953056;b=926971;opcode=110;
			#100	a=-784029;b=622893;opcode=100;
			#100	a=410076;b=-428400;opcode=001;
			#100	a=430254;b=-914116;opcode=000;
			#100	a=628362;b=-309;opcode=100;
			#100	a=-917565;b=70979;opcode=000;
			#100	a=-217247;b=280147;opcode=000;
			#100	a=157822;b=-983979;opcode=111;
			#100	a=762669;b=-258768;opcode=111;
			#100	a=993986;b=471365;opcode=001;
			#100	a=-861880;b=171502;opcode=100;
			#100	a=812861;b=-62764;opcode=000;
			#100	a=954195;b=64622;opcode=100;
			#100	a=829453;b=-958130;opcode=000;
			#100	a=279126;b=-889715;opcode=001;
			#100	a=23420;b=526879;opcode=010;
			#100	a=-349282;b=-151301;opcode=111;
			#100	a=590327;b=376101;opcode=111;
			#100	a=230426;b=-587767;opcode=110;
			#100	a=-548279;b=-137182;opcode=010;
			#100	a=395128;b=228476;opcode=001;
			#100	a=-505136;b=906577;opcode=000;
			#100	a=997851;b=917900;opcode=010;
			#100	a=651375;b=238917;opcode=110;
			#100	a=736737;b=-997081;opcode=100;
			#100	a=410544;b=621423;opcode=110;
			#100	a=654042;b=-734275;opcode=110;
			#100	a=-880561;b=601788;opcode=000;
			#100	a=-739562;b=-821980;opcode=100;
			#100	a=631254;b=820360;opcode=100;
			#100	a=68429;b=-463998;opcode=110;
			#100	a=738990;b=-695830;opcode=000;
			#100	a=262591;b=997011;opcode=111;
			#100	a=965996;b=246950;opcode=110;
			#100	a=774122;b=525862;opcode=100;
			#100	a=254082;b=-208343;opcode=010;
			#100	a=-921912;b=524409;opcode=111;
			#100	a=-570367;b=738328;opcode=010;
			#100	a=637668;b=439310;opcode=001;
			#100	a=-625304;b=-143624;opcode=110;
			#100	a=453888;b=478633;opcode=001;
			#100	a=285583;b=279888;opcode=100;
			#100	a=-284166;b=-309729;opcode=110;
			#100	a=211270;b=-617800;opcode=111;
			#100	a=627408;b=-448066;opcode=000;
			#100	a=15910;b=-546061;opcode=000;
			#100	a=-536599;b=986862;opcode=100;
			#100	a=-574701;b=568557;opcode=110;
			#100	a=705808;b=607084;opcode=100;
			#100	a=798980;b=-737225;opcode=000;
			#100	a=-200729;b=-529251;opcode=110;
			#100	a=78798;b=837754;opcode=111;
			#100	a=-94081;b=118714;opcode=010;
			#100	a=811942;b=-894060;opcode=100;
			#100	a=-166280;b=737671;opcode=100;
			#100	a=266576;b=-427176;opcode=001;
			#100	a=917673;b=-437235;opcode=010;
			#100	a=-752373;b=-646071;opcode=111;
			#100	a=-236738;b=721504;opcode=000;
			#100	a=-11710;b=-886378;opcode=110;
			#100	a=512371;b=786225;opcode=100;
			#100	a=-121576;b=-182272;opcode=001;
			#100	a=931299;b=-918227;opcode=111;
			#100	a=-103559;b=-652025;opcode=000;
			#100	a=-726491;b=500986;opcode=001;
			#100	a=75592;b=-72309;opcode=110;
			#100	a=615808;b=-495141;opcode=010;
			#100	a=-406793;b=622415;opcode=001;
			#100	a=967010;b=67446;opcode=100;
			#100	a=-607979;b=-413485;opcode=100;
			#100	a=851430;b=-148706;opcode=010;
			#100	a=778196;b=-925529;opcode=111;
			#100	a=-175018;b=-163347;opcode=001;
			#100	a=-385434;b=203071;opcode=000;
			#100	a=-472801;b=537693;opcode=111;
			#100	a=260363;b=-549761;opcode=110;
			#100	a=-230004;b=108287;opcode=010;
			#100	a=-774326;b=-474601;opcode=010;
			#100	a=-589063;b=44916;opcode=000;
			#100	a=562356;b=-788562;opcode=000;
			#100	a=551352;b=-822836;opcode=010;
			#100	a=854508;b=-629714;opcode=000;
			#100	a=331130;b=2416;opcode=100;
			#100	a=351719;b=-289040;opcode=001;
			#100	a=-334523;b=-402695;opcode=111;
			#100	a=967820;b=-607569;opcode=001;
			#100	a=-578485;b=-532482;opcode=010;
			#100	a=924802;b=-993218;opcode=010;
			#100	a=-821890;b=-991412;opcode=010;
			#100	a=829249;b=272635;opcode=110;
			#100	a=328000;b=-326138;opcode=000;
			#100	a=835980;b=562209;opcode=001;
			#100	a=-911572;b=-157258;opcode=001;
			#100	a=-605921;b=-507707;opcode=001;
			#100	a=-173242;b=-984396;opcode=010;
			#100	a=-558950;b=252079;opcode=110;
			#100	a=-187218;b=-874548;opcode=000;
			#100	a=-475335;b=-403861;opcode=111;
			#100	a=-608620;b=377328;opcode=010;
			#100	a=557753;b=-490797;opcode=010;
			#100	a=-385454;b=604052;opcode=000;
			#100	a=976481;b=191473;opcode=001;
			#100	a=933051;b=-241354;opcode=001;
			#100	a=707689;b=-750637;opcode=001;
			#100	a=-595872;b=-165417;opcode=010;
			#100	a=190602;b=-879415;opcode=110;
			#100	a=217792;b=327799;opcode=100;
			#100	a=960272;b=92422;opcode=001;
			#100	a=-294874;b=208366;opcode=000;
			#100	a=383889;b=-228080;opcode=100;
			#100	a=534091;b=-961787;opcode=110;
			#100	a=3311;b=-192;opcode=010;
			#100	a=671388;b=-289367;opcode=110;
			#100	a=357919;b=474360;opcode=100;
			#100	a=-751975;b=8898;opcode=110;
			#100	a=469607;b=117234;opcode=010;
			#100	a=495901;b=735973;opcode=110;
			#100	a=467170;b=-302485;opcode=010;
			#100	a=-90935;b=-875776;opcode=000;
			#100	a=251909;b=-252159;opcode=100;
			#100	a=463655;b=-226986;opcode=010;
			#100	a=-869175;b=-366743;opcode=000;
			#100	a=530007;b=-957112;opcode=111;
			#100	a=34200;b=174465;opcode=111;
			#100	a=300567;b=143402;opcode=000;
			#100	a=-632098;b=-812465;opcode=010;
			#100	a=-771159;b=-317095;opcode=100;
			#100	a=-193457;b=-264136;opcode=110;
			#100	a=-779022;b=94672;opcode=000;
			#100	a=459585;b=-212320;opcode=111;
			#100	a=-902230;b=506406;opcode=001;
			#100	a=-322932;b=545997;opcode=000;
			#100	a=549926;b=130807;opcode=110;
			#100	a=937446;b=841238;opcode=100;
			#100	a=884893;b=-686748;opcode=001;
			#100	a=-956285;b=-362288;opcode=100;
			#100	a=-403177;b=-932168;opcode=010;
			#100	a=335703;b=834276;opcode=110;
			#100	a=873597;b=-355342;opcode=111;
			#100	a=-523362;b=909171;opcode=111;
			#100	a=142395;b=334303;opcode=000;
			#100	a=-78921;b=242420;opcode=001;
			#100	a=-250555;b=-446779;opcode=001;
			#100	a=406976;b=831962;opcode=110;
			#100	a=878986;b=-617580;opcode=110;
			#100	a=164763;b=282902;opcode=001;
			#100	a=645336;b=206105;opcode=010;
			#100	a=873435;b=840463;opcode=010;
			#100	a=397531;b=192510;opcode=000;
			#100	a=-532681;b=-179701;opcode=111;
			#100	a=-793181;b=159132;opcode=100;
			#100	a=106532;b=959699;opcode=010;
			#100	a=-241578;b=-412944;opcode=010;
			#100	a=266265;b=611508;opcode=010;
			#100	a=-559924;b=889433;opcode=100;
			#100	a=-689802;b=-766060;opcode=110;
			#100	a=393850;b=395325;opcode=001;
			#100	a=-97650;b=400311;opcode=010;
			#100	a=-866585;b=500376;opcode=110;
			#100	a=-907198;b=-513402;opcode=000;
			#100	a=-23697;b=842302;opcode=100;
			#100	a=-102471;b=-82326;opcode=000;
			#100	a=521224;b=534897;opcode=111;
			#100	a=110356;b=770776;opcode=010;
			#100	a=50630;b=370308;opcode=001;
			#100	a=-124224;b=-9913;opcode=110;
			#100	a=-363822;b=-119382;opcode=100;
			#100	a=684381;b=355352;opcode=010;
			#100	a=185110;b=836245;opcode=111;
			#100	a=257238;b=913746;opcode=100;
			#100	a=153249;b=-396672;opcode=100;
			#100	a=-256629;b=700057;opcode=100;
			#100	a=-549597;b=-707585;opcode=100;
			#100	a=249860;b=563581;opcode=110;
			#100	a=-703958;b=-125067;opcode=110;
			#100	a=-547125;b=-72615;opcode=010;
			#100	a=928319;b=839041;opcode=100;
			#100	a=-219474;b=-453923;opcode=001;
			#100	a=-818802;b=157886;opcode=001;
			#100	a=-711432;b=922659;opcode=000;
			#100	a=622991;b=794138;opcode=100;
			#100	a=-143953;b=-813043;opcode=110;
			#100	a=665470;b=-106394;opcode=110;
			#100	a=218876;b=-156869;opcode=010;
			#100	a=115634;b=-841047;opcode=010;
			#100	a=761481;b=-776905;opcode=110;
			#100	a=-135676;b=-18893;opcode=010;
			#100	a=289882;b=-121541;opcode=001;
			#100	a=125702;b=-625282;opcode=000;
			#100	a=719859;b=461492;opcode=000;
			#100	a=-500657;b=254715;opcode=110;
			#100	a=131716;b=-611327;opcode=001;
			#100	a=441838;b=583723;opcode=000;
			#100	a=81962;b=744693;opcode=001;
			#100	a=-448386;b=490397;opcode=001;
			#100	a=635376;b=-649759;opcode=010;
			#100	a=-859338;b=-645299;opcode=010;
			#100	a=-509193;b=469276;opcode=010;
			#100	a=712033;b=255891;opcode=110;
			#100	a=514385;b=54265;opcode=111;
			#100	a=557871;b=804820;opcode=000;
			#100	a=-855388;b=-809321;opcode=111;
			#100	a=-262743;b=-710742;opcode=001;
			#100	a=911554;b=485132;opcode=110;
			#100	a=-142624;b=-669401;opcode=100;
			#100	a=519760;b=-949844;opcode=111;
			#100	a=327894;b=-576918;opcode=001;
			#100	a=-421931;b=699910;opcode=000;
			#100	a=-733982;b=-727790;opcode=100;
			#100	a=511566;b=-678908;opcode=010;
			#100	a=923044;b=74946;opcode=100;
			#100	a=143726;b=951052;opcode=010;
			#100	a=941936;b=-833080;opcode=110;
			#100	a=53694;b=150575;opcode=000;
			#100	a=160702;b=-845554;opcode=001;
			#100	a=251779;b=-727543;opcode=100;
			#100	a=-706238;b=-975144;opcode=110;
			#100	a=-121707;b=823628;opcode=110;
			#100	a=969359;b=-178621;opcode=010;
			#100	a=693790;b=-672743;opcode=111;
			#100	a=29075;b=-54884;opcode=010;
			#100	a=-667706;b=-325097;opcode=111;
			#100	a=-993333;b=-353899;opcode=000;
			#100	a=-421081;b=-650414;opcode=010;
			#100	a=909186;b=20977;opcode=000;
			#100	a=249251;b=-226717;opcode=100;
			#100	a=928119;b=-11221;opcode=111;
			#100	a=-235628;b=848190;opcode=001;
			#100	a=-79374;b=943943;opcode=110;
			#100	a=970330;b=483446;opcode=110;
			#100	a=433914;b=-766822;opcode=000;
			#100	a=221394;b=616665;opcode=110;
			#100	a=-307426;b=-569430;opcode=110;
			#100	a=125635;b=134029;opcode=100;
			#100	a=732499;b=-871617;opcode=010;
			#100	a=978980;b=652963;opcode=000;
			#100	a=-751169;b=996578;opcode=100;
			#100	a=-797043;b=615955;opcode=001;
			#100	a=332038;b=-856150;opcode=110;
			#100	a=-584308;b=-93185;opcode=111;
			#100	a=21805;b=-385071;opcode=111;
			#100	a=139909;b=519761;opcode=001;
			#100	a=838920;b=-671171;opcode=010;
			#100	a=870449;b=-169130;opcode=001;
			#100	a=-992544;b=-501325;opcode=100;
			#100	a=-494518;b=-468141;opcode=010;
			#100	a=593899;b=-269071;opcode=100;
			#100	a=-747333;b=835939;opcode=000;
			#100	a=-207291;b=288821;opcode=100;
			#100	a=-697011;b=620399;opcode=111;
			#100	a=763826;b=-48024;opcode=100;
			#100	a=-161463;b=324165;opcode=010;
			#100	a=564461;b=-70023;opcode=110;
			#100	a=-179307;b=624330;opcode=111;
			#100	a=-420310;b=-372256;opcode=010;
			#100	a=390474;b=-341833;opcode=111;
			#100	a=-861134;b=80053;opcode=000;
			#100	a=722030;b=239645;opcode=001;
			#100	a=-967275;b=519646;opcode=111;
			#100	a=167469;b=692588;opcode=001;
			#100	a=-608602;b=224972;opcode=100;
			#100	a=828545;b=930792;opcode=010;
			#100	a=362130;b=24924;opcode=000;
			#100	a=-187928;b=324058;opcode=010;
			#100	a=165385;b=-718329;opcode=010;
			#100	a=-236795;b=-835677;opcode=110;
			#100	a=364419;b=-82754;opcode=110;
			#100	a=-106107;b=-636634;opcode=110;
			#100	a=-516600;b=-502623;opcode=000;
			#100	a=904119;b=639549;opcode=001;
			#100	a=-118384;b=-570063;opcode=111;
			#100	a=-87299;b=227667;opcode=010;
			#100	a=247371;b=-954691;opcode=111;
			#100	a=186063;b=-8517;opcode=010;
			#100	a=115816;b=-854450;opcode=111;
			#100	a=20259;b=219304;opcode=100;
			#100	a=327991;b=-871315;opcode=010;
			#100	a=861396;b=186917;opcode=100;
			#100	a=-378603;b=-360679;opcode=001;
			#100	a=-426247;b=305081;opcode=001;
			#100	a=431317;b=692158;opcode=001;
			#100	a=553875;b=-353461;opcode=100;
			#100	a=128219;b=360969;opcode=100;
			#100	a=789885;b=-684220;opcode=010;
			#100	a=-330566;b=283873;opcode=001;
			#100	a=301237;b=297810;opcode=010;
			#100	a=-338750;b=23486;opcode=010;
			#100	a=-927860;b=-203068;opcode=110;
			#100	a=334360;b=29490;opcode=001;
			#100	a=717877;b=625799;opcode=001;
			#100	a=-177897;b=-828477;opcode=010;
			#100	a=812216;b=-122477;opcode=000;
			#100	a=555040;b=917311;opcode=000;
			#100	a=-98616;b=-939304;opcode=010;
			#100	a=359220;b=-988853;opcode=000;
			#100	a=542700;b=53701;opcode=000;
			#100	a=-338774;b=-795213;opcode=110;
			#100	a=-955403;b=-418850;opcode=001;
			#100	a=458345;b=887047;opcode=110;
			#100	a=-368027;b=818259;opcode=000;
			#100	a=-349117;b=628734;opcode=000;
			#100	a=-646801;b=-466152;opcode=001;
			#100	a=733259;b=-903676;opcode=000;
			#100	a=249494;b=532992;opcode=100;
			#100	a=921114;b=936044;opcode=001;
			#100	a=592156;b=774785;opcode=000;
			#100	a=445509;b=-879913;opcode=001;
			#100	a=-423587;b=-244245;opcode=010;
			#100	a=52442;b=335809;opcode=111;
			#100	a=-266823;b=569571;opcode=010;
			#100	a=765223;b=-478202;opcode=001;
			#100	a=948610;b=-132254;opcode=110;
			#100	a=-488246;b=-243071;opcode=010;
			#100	a=-826125;b=-787044;opcode=111;
			#100	a=-601792;b=-570320;opcode=001;
			#100	a=-64768;b=209225;opcode=000;
			#100	a=490754;b=604716;opcode=110;
			#100	a=542620;b=-172647;opcode=010;
			#100	a=185003;b=-895329;opcode=000;
			#100	a=39595;b=876565;opcode=010;
			#100	a=-650582;b=-897087;opcode=110;
			#100	a=269850;b=812097;opcode=111;
			#100	a=589137;b=-578951;opcode=001;
			#100	a=-918807;b=314112;opcode=010;
			#100	a=-918466;b=144766;opcode=111;
			#100	a=241285;b=-423744;opcode=010;
			#100	a=-718579;b=570701;opcode=100;
			#100	a=513124;b=-828467;opcode=010;
			#100	a=-905951;b=19145;opcode=100;
			#100	a=2636;b=-691406;opcode=001;
			#100	a=-422680;b=-994645;opcode=001;
			#100	a=113389;b=-395908;opcode=000;
			#100	a=-169303;b=-232360;opcode=001;
			#100	a=-283711;b=-256734;opcode=110;
			#100	a=706896;b=-578388;opcode=100;
			#100	a=595087;b=-736137;opcode=000;
			#100	a=-84167;b=-921685;opcode=100;
			#100	a=-224803;b=108034;opcode=010;
			#100	a=564676;b=357066;opcode=000;
			#100	a=-435712;b=-819696;opcode=001;
			#100	a=773800;b=-575936;opcode=111;
			#100	a=-950449;b=62922;opcode=111;
			#100	a=514443;b=201263;opcode=010;
			#100	a=-170528;b=838230;opcode=010;
			#100	a=428293;b=553319;opcode=001;
			#100	a=-628047;b=709474;opcode=100;
			#100	a=-425021;b=295620;opcode=110;
			#100	a=-143047;b=-474014;opcode=100;
			#100	a=200647;b=25983;opcode=010;
			#100	a=411834;b=-184347;opcode=000;
			#100	a=-589391;b=525734;opcode=110;
			#100	a=-889558;b=41836;opcode=000;
			#100	a=22611;b=-785403;opcode=000;
			#100	a=129646;b=598856;opcode=110;
			#100	a=177566;b=-910241;opcode=111;
			#100	a=-515585;b=-409182;opcode=001;
			#100	a=776799;b=669683;opcode=000;
			#100	a=-280796;b=-228769;opcode=000;
			#100	a=654541;b=189954;opcode=111;
			#100	a=-243119;b=244305;opcode=000;
			#100	a=-504754;b=-78526;opcode=110;
			#100	a=201236;b=758596;opcode=111;
			#100	a=-517407;b=-70654;opcode=100;
			#100	a=440198;b=-616500;opcode=000;
			#100	a=-263497;b=-639589;opcode=111;
			#100	a=-556007;b=-309571;opcode=111;
			#100	a=114296;b=-818749;opcode=010;
			#100	a=-790207;b=-319097;opcode=000;
			#100	a=-262262;b=-502299;opcode=110;
			#100	a=-840137;b=345150;opcode=111;
			#100	a=-807003;b=122074;opcode=111;
			#100	a=730043;b=-211435;opcode=111;
			#100	a=-177575;b=-867744;opcode=000;
			#100	a=-293174;b=696935;opcode=111;
			#100	a=944420;b=-492537;opcode=010;
			#100	a=-343987;b=-57063;opcode=001;
			#100	a=-730307;b=155133;opcode=000;
			#100	a=337759;b=386187;opcode=010;
			#100	a=-287176;b=-469375;opcode=111;
			#100	a=-401195;b=-398713;opcode=001;
			#100	a=-673277;b=-245852;opcode=010;
			#100	a=-740148;b=-630008;opcode=001;
			#100	a=-67783;b=-576648;opcode=000;
			#100	a=11782;b=-569290;opcode=010;
			#100	a=598104;b=-597362;opcode=110;
			#100	a=954102;b=715802;opcode=000;
			#100	a=776782;b=-59891;opcode=100;
			#100	a=-353525;b=375849;opcode=000;
			#100	a=-23063;b=-327071;opcode=010;
			#100	a=992221;b=211337;opcode=110;
			#100	a=581805;b=-558373;opcode=100;
			#100	a=367767;b=-682823;opcode=010;
			#100	a=-597050;b=-682712;opcode=110;
			#100	a=-492268;b=-804576;opcode=100;
			#100	a=-698961;b=-9312;opcode=100;
			#100	a=351146;b=-691019;opcode=001;
			#100	a=559021;b=602674;opcode=000;
			#100	a=-17032;b=-557736;opcode=010;
			#100	a=85012;b=551208;opcode=010;
			#100	a=-76265;b=-831465;opcode=000;
			#100	a=897930;b=894987;opcode=100;
			#100	a=13548;b=551407;opcode=001;
			#100	a=98460;b=244971;opcode=001;
			#100	a=792472;b=481936;opcode=100;
			#100	a=-157682;b=-572321;opcode=111;
			#100	a=-522072;b=-721988;opcode=110;
			#100	a=-120409;b=-408373;opcode=000;
			#100	a=-996699;b=-648581;opcode=100;
			#100	a=658047;b=116454;opcode=111;
			#100	a=-260724;b=-362443;opcode=111;
			#100	a=-198214;b=-273532;opcode=001;
			#100	a=-985706;b=955974;opcode=111;
			#100	a=-870676;b=626228;opcode=111;
			#100	a=929916;b=830141;opcode=110;
			#100	a=-496132;b=556600;opcode=110;
			#100	a=-518340;b=599072;opcode=111;
			#100	a=-176336;b=582719;opcode=001;
			#100	a=467351;b=-843269;opcode=001;
			#100	a=729592;b=-746630;opcode=110;
			#100	a=-585765;b=986578;opcode=100;
			#100	a=617669;b=388222;opcode=001;
			#100	a=821132;b=990013;opcode=001;
			#100	a=272172;b=723222;opcode=001;
			#100	a=143677;b=-618329;opcode=000;
			#100	a=859415;b=59098;opcode=000;
			#100	a=-989101;b=901052;opcode=111;
			#100	a=-913987;b=94944;opcode=001;
			#100	a=-580807;b=791096;opcode=110;
			#100	a=-408154;b=425670;opcode=000;
			#100	a=41765;b=74211;opcode=111;
			#100	a=817920;b=758102;opcode=000;
			#100	a=-244221;b=777615;opcode=010;
			#100	a=-728796;b=757972;opcode=100;
			#100	a=735051;b=1309;opcode=000;
			#100	a=416508;b=664488;opcode=100;
			#100	a=358181;b=920257;opcode=100;
			#100	a=771890;b=949426;opcode=010;
			#100	a=-689035;b=818886;opcode=111;
			#100	a=-576304;b=-273452;opcode=110;
			#100	a=-596749;b=-269300;opcode=111;
			#100	a=-958869;b=201830;opcode=000;
			#100	a=823127;b=-670184;opcode=001;
			#100	a=-296812;b=354414;opcode=111;
			#100	a=345290;b=-87490;opcode=111;
			#100	a=168920;b=32568;opcode=111;
			#100	a=-852578;b=-202811;opcode=100;
			#100	a=-753497;b=670876;opcode=010;
			#100	a=636296;b=384589;opcode=100;
			#100	a=972431;b=-85701;opcode=010;
			#100	a=621881;b=446375;opcode=100;
			#100	a=-302108;b=-793258;opcode=111;
			#100	a=923694;b=-177248;opcode=000;
			#100	a=-403704;b=831399;opcode=111;
			#100	a=185941;b=681870;opcode=001;
			#100	a=-749863;b=-611568;opcode=110;
			#100	a=936317;b=-68664;opcode=001;
			#100	a=-891482;b=37925;opcode=100;
			#100	a=315224;b=-723958;opcode=001;
			#100	a=949989;b=-570237;opcode=010;
			#100	a=-353576;b=-49284;opcode=100;
			#100	a=-15312;b=-207934;opcode=100;
			#100	a=-152770;b=404602;opcode=001;
			#100	a=706743;b=-842303;opcode=001;
			#100	a=-29027;b=455221;opcode=010;
			#100	a=-954054;b=153631;opcode=010;
			#100	a=131611;b=-452901;opcode=110;
			#100	a=68682;b=-463755;opcode=110;
			#100	a=-375438;b=558540;opcode=001;
			#100	a=-915516;b=-287120;opcode=111;
			#100	a=536530;b=603166;opcode=001;
			#100	a=831137;b=-795648;opcode=110;
			#100	a=-36751;b=234264;opcode=010;
			#100	a=-232384;b=43365;opcode=010;
			#100	a=-160279;b=964863;opcode=000;
			#100	a=960183;b=-637506;opcode=111;
			#100	a=217631;b=660391;opcode=000;
			#100	a=-985548;b=-293305;opcode=010;
			#100	a=-128891;b=975772;opcode=111;
			#100	a=916729;b=-248105;opcode=000;
			#100	a=-856187;b=-918753;opcode=100;
			#100	a=-966908;b=151105;opcode=001;
			#100	a=-810681;b=174172;opcode=001;
			#100	a=-676011;b=-241090;opcode=001;
			#100	a=-742850;b=-375434;opcode=100;
			#100	a=-347117;b=-275908;opcode=111;
			#100	a=-972946;b=537392;opcode=100;
			#100	a=-435932;b=351372;opcode=001;
			#100	a=880397;b=-363146;opcode=100;
			#100	a=-242991;b=506308;opcode=100;
			#100	a=-287665;b=360614;opcode=100;
			#100	a=146549;b=336896;opcode=100;
			#100	a=-39132;b=59310;opcode=001;
			#100	a=-894141;b=-800977;opcode=000;
			#100	a=-90188;b=-564099;opcode=111;
			#100	a=-458539;b=-627614;opcode=000;
			#100	a=-309001;b=-71858;opcode=111;
			#100	a=-136372;b=561349;opcode=000;
			#100	a=455745;b=557380;opcode=110;
			#100	a=-111941;b=-821366;opcode=010;
			#100	a=-602061;b=-430422;opcode=001;
			#100	a=946917;b=354958;opcode=001;
			#100	a=568467;b=894751;opcode=111;
			#100	a=192625;b=-785406;opcode=111;
			#100	a=928948;b=163461;opcode=110;
			#100	a=-625779;b=-319698;opcode=111;
			#100	a=692218;b=455122;opcode=111;
			#100	a=606549;b=-400612;opcode=111;
			#100	a=-940623;b=-70137;opcode=110;
			#100	a=340518;b=-466575;opcode=111;
			#100	a=-530640;b=38497;opcode=000;
			#100	a=180059;b=611498;opcode=100;
			#100	a=8240;b=680950;opcode=111;
			#100	a=665056;b=-524555;opcode=000;
			#100	a=-199398;b=240452;opcode=000;
			#100	a=-898610;b=154506;opcode=010;
			#100	a=-342555;b=405807;opcode=100;
			#100	a=-853741;b=-414793;opcode=010;
			#100	a=158321;b=225910;opcode=000;
			#100	a=236934;b=28406;opcode=000;
			#100	a=822444;b=875130;opcode=010;
			#100	a=-103864;b=203372;opcode=010;
			#100	a=-119881;b=-852300;opcode=010;
			#100	a=-280576;b=-928174;opcode=001;
			#100	a=-215167;b=-542202;opcode=010;
			#100	a=-612286;b=502907;opcode=001;
			#100	a=756290;b=-552740;opcode=110;
			#100	a=824099;b=908671;opcode=110;
			#100	a=229095;b=-22619;opcode=000;
			#100	a=571505;b=-376870;opcode=000;
			#100	a=-739317;b=14346;opcode=001;
			#100	a=142935;b=913359;opcode=110;
			#100	a=467583;b=-379879;opcode=111;
			#100	a=-839352;b=903658;opcode=100;
			#100	a=108783;b=-440847;opcode=111;
			#100	a=213673;b=-133308;opcode=001;
			#100	a=629280;b=-892290;opcode=000;
			#100	a=-822230;b=-511958;opcode=111;
			#100	a=-35747;b=932102;opcode=100;
			#100	a=691147;b=422777;opcode=010;
			#100	a=-251879;b=566776;opcode=100;
			#100	a=511274;b=-806431;opcode=001;
			#100	a=362243;b=957894;opcode=111;
			#100	a=280785;b=589628;opcode=111;
			#100	a=-92695;b=677702;opcode=000;
			#100	a=634891;b=298865;opcode=111;
			#100	a=-15088;b=-424341;opcode=001;
			#100	a=-712445;b=-456030;opcode=100;
			#100	a=-532635;b=922260;opcode=010;
			#100	a=-988630;b=-17926;opcode=010;
			#100	a=-865388;b=349412;opcode=010;
			#100	a=222104;b=266328;opcode=010;
			#100	a=786712;b=-745161;opcode=110;
			#100	a=-822159;b=723376;opcode=110;
			#100	a=439918;b=-364496;opcode=010;
			#100	a=718605;b=570181;opcode=010;
			#100	a=947313;b=-890955;opcode=010;
			#100	a=878658;b=948380;opcode=110;
			#100	a=-833337;b=-744862;opcode=001;
			#100	a=774430;b=627366;opcode=001;
			#100	a=222230;b=-54372;opcode=111;
			#100	a=-270312;b=381642;opcode=000;
			#100	a=-961823;b=-995061;opcode=100;
			#100	a=-726153;b=-241165;opcode=110;
			#100	a=-240858;b=-202573;opcode=100;
			#100	a=790327;b=-40740;opcode=111;
			#100	a=-613075;b=-471283;opcode=010;
			#100	a=-698811;b=-831664;opcode=100;
			#100	a=-890523;b=876398;opcode=000;
			#100	a=-979801;b=495760;opcode=001;
			#100	a=-543672;b=-615862;opcode=001;
			#100	a=-707614;b=-969316;opcode=111;
			#100	a=-592242;b=-970128;opcode=010;
			#100	a=-289067;b=858443;opcode=001;
			#100	a=-351055;b=755763;opcode=100;
			#100	a=546618;b=208983;opcode=000;
			#100	a=-264433;b=28624;opcode=111;
			#100	a=155461;b=-979531;opcode=110;
			#100	a=-329418;b=900963;opcode=100;
			#100	a=-653745;b=630401;opcode=001;
			#100	a=-483604;b=-482932;opcode=000;
			#100	a=305341;b=-166365;opcode=110;
			#100	a=-580452;b=-331139;opcode=100;
			#100	a=303744;b=362515;opcode=000;
			#100	a=-143552;b=-981435;opcode=000;
			#100	a=-392020;b=-313020;opcode=110;
			#100	a=-120355;b=-461150;opcode=110;
			#100	a=250861;b=-353644;opcode=001;
			#100	a=-128981;b=418861;opcode=111;
			#100	a=230641;b=-277682;opcode=110;
			#100	a=-953905;b=-67545;opcode=001;
			#100	a=970852;b=130112;opcode=001;
			#100	a=345231;b=780408;opcode=110;
			#100	a=-849155;b=363732;opcode=001;
			#100	a=38670;b=-948486;opcode=110;
			#100	a=-178609;b=171585;opcode=111;
			#100	a=-956518;b=-775846;opcode=000;
			#100	a=473014;b=-688817;opcode=010;
			#100	a=330000;b=100348;opcode=110;
			#100	a=626623;b=18752;opcode=000;
			#100	a=-995393;b=457107;opcode=000;
			#100	a=290402;b=238753;opcode=100;
			#100	a=349450;b=864121;opcode=001;
			#100	a=-303465;b=-559924;opcode=010;
			#100	a=357621;b=-23974;opcode=110;
			#100	a=-310423;b=-161270;opcode=100;
			#100	a=-552950;b=-95642;opcode=001;
			#100	a=179152;b=231667;opcode=100;
			#100	a=-713948;b=-371677;opcode=001;
			#100	a=-238363;b=242860;opcode=111;
			#100	a=92103;b=-387927;opcode=111;
			#100	a=630529;b=-420523;opcode=111;
			#100	a=858026;b=790825;opcode=110;
			#100	a=-928224;b=361021;opcode=000;
			#100	a=-922405;b=-330837;opcode=110;
			#100	a=-839205;b=27705;opcode=000;
			#100	a=232284;b=413508;opcode=001;
			#100	a=139205;b=908531;opcode=000;
			#100	a=-231363;b=565955;opcode=100;
			#100	a=432093;b=358841;opcode=111;
			#100	a=-168355;b=532408;opcode=110;
			#100	a=745796;b=214283;opcode=110;
			#100	a=-381039;b=306844;opcode=111;
			#100	a=-82873;b=954017;opcode=111;
			#100	a=-371694;b=-780404;opcode=100;
			#100	a=-849350;b=1544;opcode=100;
			#100	a=466405;b=-672021;opcode=001;
			#100	a=430032;b=-673972;opcode=001;
			#100	a=567275;b=-641844;opcode=001;
			#100	a=-341150;b=514098;opcode=010;
			#100	a=-103095;b=-613339;opcode=111;
			#100	a=935013;b=566627;opcode=001;
			#100	a=-395483;b=779565;opcode=000;
			#100	a=-750884;b=-573014;opcode=001;
			#100	a=-185277;b=-586691;opcode=000;
			#100	a=355041;b=15130;opcode=110;
			#100	a=-393894;b=684403;opcode=001;
			#100	a=-299941;b=-365834;opcode=001;
			#100	a=-485208;b=-700233;opcode=100;
			#100	a=-944497;b=-694616;opcode=000;
			#100	a=-906359;b=-141299;opcode=001;
			#100	a=-485984;b=509121;opcode=000;
			#100	a=-351337;b=-500345;opcode=000;
			#100	a=-311563;b=-892139;opcode=100;
			#100	a=324616;b=671957;opcode=100;
			#100	a=-573255;b=-186115;opcode=100;
			#100	a=561160;b=-245041;opcode=010;
			#100	a=-999023;b=328721;opcode=000;
			#100	a=-391597;b=-21686;opcode=100;
			#100	a=939936;b=698919;opcode=111;
			#100	a=424087;b=-50019;opcode=110;
			#100	a=-731542;b=-950592;opcode=100;
			#100	a=651166;b=-943730;opcode=100;
			#100	a=208153;b=-813432;opcode=100;
			#100	a=684029;b=302610;opcode=111;
			#100	a=199656;b=-344876;opcode=110;
			#100	a=-353940;b=953990;opcode=110;
			#100	a=-722666;b=786939;opcode=110;
			#100	a=-45107;b=-396524;opcode=111;
			#100	a=-747463;b=995934;opcode=001;
			#100	a=488582;b=520687;opcode=001;
			#100	a=-691769;b=468295;opcode=001;
			#100	a=-775118;b=-488868;opcode=111;
			#100	a=657546;b=-197820;opcode=100;
			#100	a=-475445;b=-138834;opcode=111;
			#100	a=209866;b=259257;opcode=001;
			#100	a=370689;b=-287694;opcode=001;
			#100	a=99000;b=-194159;opcode=010;
			#100	a=906826;b=-468131;opcode=110;
			#100	a=-611039;b=-380628;opcode=110;
			#100	a=-500115;b=-862313;opcode=100;
			#100	a=872185;b=83796;opcode=110;
			#100	a=779803;b=266295;opcode=100;
			#100	a=894322;b=298884;opcode=100;
			#100	a=-716423;b=-172772;opcode=111;
			#100	a=-533517;b=244920;opcode=100;
			#100	a=-572286;b=-558738;opcode=111;
			#100	a=374025;b=-825224;opcode=010;
			#100	a=495878;b=-358361;opcode=111;
			#100	a=143930;b=212718;opcode=100;
			#100	a=710084;b=-886880;opcode=001;
			#100	a=-114907;b=-830638;opcode=111;
			#100	a=-858766;b=298739;opcode=001;
			#100	a=732325;b=-204098;opcode=100;
			#100	a=851407;b=103745;opcode=010;
			#100	a=-174049;b=-653994;opcode=111;
			#100	a=-303292;b=447512;opcode=110;
			#100	a=-242154;b=-816075;opcode=111;
			#100	a=-276080;b=-476912;opcode=010;
			#100	a=126974;b=-743324;opcode=100;
			#100	a=-478381;b=-451304;opcode=110;
			#100	a=-121512;b=759107;opcode=111;
			#100	a=-947905;b=115823;opcode=100;
			#100	a=-207015;b=714935;opcode=001;
			#100	a=-495711;b=-325862;opcode=001;
			#100	a=-835471;b=192149;opcode=100;
			#100	a=-116872;b=-38551;opcode=110;
			#100	a=-573695;b=883778;opcode=001;
			#100	a=-877598;b=672983;opcode=110;
			#100	a=742430;b=-501525;opcode=110;
			#100	a=736209;b=-575585;opcode=001;
			#100	a=-550650;b=-462062;opcode=000;
			#100	a=286014;b=-76885;opcode=110;
			#100	a=261587;b=906916;opcode=111;
			#100	a=916539;b=373224;opcode=111;
			#100	a=266685;b=-187822;opcode=010;
			#100	a=233746;b=78146;opcode=000;
			#100	a=-271387;b=202783;opcode=100;
			#100	a=-273694;b=-46902;opcode=000;
			#100	a=-592095;b=-743747;opcode=010;
			#100	a=402335;b=-486499;opcode=010;
			#100	a=867055;b=471814;opcode=110;
			#100	a=446451;b=784822;opcode=000;
			#100	a=-198193;b=-426277;opcode=000;
			#100	a=-130125;b=-482928;opcode=010;
			#100	a=-446313;b=-353431;opcode=000;
			#100	a=-627988;b=570687;opcode=001;
			#100	a=711493;b=-902028;opcode=001;
			#100	a=-983296;b=-413147;opcode=110;
			#100	a=280036;b=-736245;opcode=010;
			#100	a=151454;b=-27064;opcode=010;
			#100	a=620918;b=968110;opcode=010;
			#100	a=-330749;b=504033;opcode=100;
			#100	a=-721310;b=333172;opcode=111;
			#100	a=-755551;b=462771;opcode=001;
			#100	a=-895697;b=-71849;opcode=100;
			#100	a=57755;b=-30600;opcode=110;
			#100	a=-975765;b=638481;opcode=010;
			#100	a=612955;b=830051;opcode=110;
			#100	a=-47016;b=-498326;opcode=110;
			#100	a=-533944;b=511457;opcode=010;
			#100	a=-328479;b=-763313;opcode=001;
			#100	a=-296497;b=360215;opcode=001;
			#100	a=888362;b=115316;opcode=100;
			#100	a=-758697;b=984056;opcode=100;
			#100	a=-860377;b=-910533;opcode=100;
			#100	a=310250;b=-322584;opcode=000;
			#100	a=-976271;b=110900;opcode=100;
			#100	a=967503;b=719503;opcode=010;
			#100	a=-993205;b=-731438;opcode=010;
			#100	a=539461;b=-93357;opcode=010;
			#100	a=945481;b=-891548;opcode=100;
			#100	a=-666943;b=398065;opcode=001;
			#100	a=-390583;b=802199;opcode=110;
			#100	a=-289855;b=824477;opcode=100;
			#100	a=-871825;b=464004;opcode=111;
			#100	a=186593;b=-516369;opcode=111;
			#100	a=100592;b=69303;opcode=001;
			#100	a=911925;b=-188170;opcode=110;
			#100	a=731178;b=17012;opcode=010;
			#100	a=970616;b=-583981;opcode=110;
			#100	a=-782254;b=57543;opcode=010;
			#100	a=631860;b=8757;opcode=000;
			#100	a=636075;b=377371;opcode=100;
			#100	a=-964543;b=732702;opcode=110;
			#100	a=444143;b=-8240;opcode=010;
			#100	a=-705297;b=608265;opcode=000;
			#100	a=547819;b=-617322;opcode=010;
			#100	a=-257041;b=-804115;opcode=010;
			#100	a=-623072;b=68383;opcode=110;
			#100	a=626998;b=973192;opcode=111;
			#100	a=652136;b=-390829;opcode=110;
			#100	a=-226687;b=-89216;opcode=110;
			#100	a=-462567;b=617912;opcode=010;
			#100	a=-265366;b=-888439;opcode=001;
			#100	a=731149;b=706369;opcode=100;
			#100	a=-258875;b=305658;opcode=111;
			#100	a=-564950;b=238006;opcode=001;
			#100	a=723086;b=288430;opcode=111;
			#100	a=-18862;b=355700;opcode=000;
			#100	a=-71158;b=363776;opcode=000;
			#100	a=-249375;b=-118392;opcode=111;
			#100	a=904065;b=-228419;opcode=110;
			#100	a=-608253;b=-48812;opcode=111;
			#100	a=-499619;b=-229172;opcode=110;
			#100	a=719054;b=-569766;opcode=111;
			#100	a=-305879;b=693440;opcode=111;
			#100	a=-846591;b=-355361;opcode=010;
			#100	a=634506;b=437550;opcode=110;
			#100	a=-807335;b=-661742;opcode=110;
			#100	a=-287955;b=-448110;opcode=001;
			#100	a=-692255;b=770428;opcode=100;
			#100	a=883844;b=-392827;opcode=110;
			#100	a=985952;b=-374508;opcode=010;
			#100	a=213851;b=-857801;opcode=001;
			#100	a=-653683;b=248715;opcode=110;
			#100	a=-275505;b=-625012;opcode=001;
			#100	a=-286001;b=-542143;opcode=010;
			#100	a=-544526;b=719949;opcode=110;
			#100	a=269861;b=325507;opcode=010;
			#100	a=-259218;b=387488;opcode=000;
			#100	a=-269404;b=504687;opcode=010;
			#100	a=-402996;b=148920;opcode=100;
			#100	a=-729977;b=300676;opcode=100;
			#100	a=861973;b=545802;opcode=010;
			#100	a=-616798;b=788596;opcode=001;
			#100	a=-148744;b=-592678;opcode=110;
			#100	a=-94046;b=329199;opcode=110;
			#100	a=299601;b=142560;opcode=111;
			#100	a=399239;b=296731;opcode=000;
			#100	a=493434;b=-207578;opcode=100;
			#100	a=145072;b=405902;opcode=110;
			#100	a=-327084;b=437491;opcode=010;
			#100	a=793478;b=-852268;opcode=001;
			#100	a=-111232;b=-106779;opcode=010;
			#100	a=-13843;b=-943576;opcode=100;
			#100	a=120145;b=-132192;opcode=111;
			#100	a=141370;b=-752952;opcode=001;
			#100	a=852618;b=-692286;opcode=111;
			#100	a=-244500;b=-983553;opcode=000;
			#100	a=996237;b=721174;opcode=010;
			#100	a=-844127;b=451626;opcode=010;
			#100	a=-389943;b=-928264;opcode=001;
			#100	a=-356508;b=-514769;opcode=110;
			#100	a=894171;b=-993744;opcode=110;
			#100	a=-334800;b=-886638;opcode=000;
			#100	a=-696942;b=-842099;opcode=110;
			#100	a=-228879;b=498233;opcode=110;
			#100	a=146404;b=-285357;opcode=111;
			#100	a=-563100;b=96518;opcode=000;
			#100	a=766861;b=-414528;opcode=010;
			#100	a=-525509;b=-143040;opcode=100;
			#100	a=972141;b=270287;opcode=000;
			#100	a=-96371;b=253172;opcode=010;
			#100	a=-54551;b=-47249;opcode=111;
			#100	a=917522;b=-583889;opcode=001;
			#100	a=535637;b=-413057;opcode=000;
			#100	a=-7232;b=-213046;opcode=001;
			#100	a=410127;b=-762854;opcode=110;
			#100	a=-672333;b=-590235;opcode=111;
			#100	a=-202974;b=-634276;opcode=110;
			#100	a=503731;b=-851897;opcode=010;
			#100	a=757850;b=-570889;opcode=000;
			#100	a=-542527;b=988665;opcode=001;
			#100	a=-896164;b=160130;opcode=110;
			#100	a=409278;b=-621377;opcode=111;
			#100	a=-531093;b=443273;opcode=000;
			#100	a=317963;b=695060;opcode=100;
			#100	a=-406446;b=-663697;opcode=010;
			#100	a=-215564;b=818212;opcode=001;
			#100	a=735350;b=631018;opcode=111;
			#100	a=348453;b=830354;opcode=001;
			#100	a=461597;b=891049;opcode=111;
			#100	a=49929;b=755413;opcode=001;
			#100	a=-211904;b=746815;opcode=100;
			#100	a=-524026;b=-821671;opcode=110;
			#100	a=971886;b=-373098;opcode=001;
			#100	a=253131;b=-998789;opcode=111;
			#100	a=-14417;b=-920079;opcode=100;
			#100	a=-859613;b=988438;opcode=000;
			#100	a=-113484;b=-397321;opcode=100;
			#100	a=162018;b=-346896;opcode=110;
			#100	a=624298;b=-254853;opcode=111;
			#100	a=421667;b=576130;opcode=100;
			#100	a=618050;b=-483187;opcode=111;
			#100	a=-40332;b=-12220;opcode=100;
			#100	a=-698463;b=925280;opcode=110;
			#100	a=-62795;b=641813;opcode=110;
			#100	a=694416;b=-175293;opcode=001;
			#100	a=-145287;b=888256;opcode=100;
			#100	a=681360;b=-449367;opcode=001;
			#100	a=-952824;b=-554444;opcode=001;
			#100	a=241548;b=587600;opcode=001;
			#100	a=379018;b=-839525;opcode=111;
			#100	a=-280725;b=716692;opcode=100;
			#100	a=852287;b=533254;opcode=010;
			#100	a=-139209;b=751633;opcode=111;
			#100	a=-297248;b=-844499;opcode=100;
			#100	a=809955;b=684094;opcode=000;
			#100	a=-642635;b=147168;opcode=100;
			#100	a=-152115;b=-26354;opcode=111;
			#100	a=-201107;b=384051;opcode=110;
			#100	a=-929230;b=685360;opcode=000;
			#100	a=-912451;b=944256;opcode=111;
			#100	a=731560;b=948136;opcode=111;
			#100	a=-818913;b=593419;opcode=010;
			#100	a=-207799;b=-87560;opcode=111;
			#100	a=-849671;b=291856;opcode=111;
			#100	a=27123;b=-888004;opcode=001;
			#100	a=572857;b=-415785;opcode=111;
			#100	a=398868;b=-658844;opcode=111;
			#100	a=266102;b=976379;opcode=010;
			#100	a=645294;b=-445457;opcode=111;
			#100	a=-972605;b=-329682;opcode=010;
			#100	a=-215829;b=-663898;opcode=110;
			#100	a=824266;b=-127930;opcode=000;
			#100	a=-976842;b=-555943;opcode=100;
			#100	a=-563940;b=626123;opcode=100;
			#100	a=476675;b=394771;opcode=111;
			#100	a=-326913;b=223042;opcode=000;
			#100	a=640256;b=829301;opcode=110;
			#100	a=-61922;b=88911;opcode=000;
			#100	a=-947428;b=890810;opcode=111;
			#100	a=-431897;b=836712;opcode=001;
			#100	a=-610363;b=-832958;opcode=000;
			#100	a=529526;b=-406784;opcode=100;
			#100	a=-95691;b=-696791;opcode=110;
			#100	a=-586038;b=-776474;opcode=110;
			#100	a=-786995;b=312792;opcode=000;
			#100	a=-662923;b=-30870;opcode=001;
			#100	a=-947974;b=-365151;opcode=000;
			#100	a=852224;b=-417260;opcode=010;
			#100	a=599726;b=783314;opcode=111;
			#100	a=507487;b=-721816;opcode=110;
			#100	a=864436;b=-24742;opcode=111;
			#100	a=-512769;b=877793;opcode=001;
			#100	a=-899825;b=-561148;opcode=010;
			#100	a=-630903;b=-668033;opcode=010;
			#100	a=-789981;b=-816353;opcode=111;
			#100	a=-834359;b=-357766;opcode=100;
			#100	a=-882974;b=-167800;opcode=001;
			#100	a=-362951;b=-151305;opcode=100;
			#100	a=515528;b=-718423;opcode=000;
			#100	a=-828565;b=-770605;opcode=010;
			#100	a=597779;b=-365000;opcode=110;
			#100	a=68018;b=902058;opcode=111;
			#100	a=275892;b=347938;opcode=000;
			#100	a=-392013;b=506008;opcode=001;
			#100	a=280371;b=102023;opcode=010;
			#100	a=531483;b=802418;opcode=001;
			#100	a=912823;b=-225072;opcode=110;
			#100	a=-779917;b=93137;opcode=001;
			#100	a=196631;b=952233;opcode=110;
			#100	a=-956856;b=129350;opcode=001;
			#100	a=872736;b=63041;opcode=111;
			#100	a=-148216;b=563207;opcode=100;
			#100	a=-174468;b=-590531;opcode=111;
			#100	a=873860;b=576042;opcode=001;
			#100	a=-989811;b=-629615;opcode=111;
			#100	a=-840323;b=651085;opcode=010;
			#100	a=-877015;b=-328254;opcode=010;
			#100	a=-690038;b=-639910;opcode=110;
			#100	a=915956;b=93901;opcode=111;
			#100	a=-752504;b=-244230;opcode=100;
			#100	a=96831;b=243192;opcode=110;
			#100	a=-268238;b=-945172;opcode=111;
			#100	a=986262;b=119132;opcode=000;
			#100	a=-704198;b=675464;opcode=000;
			#100	a=-218693;b=386286;opcode=001;
			#100	a=-958555;b=35120;opcode=010;
			#100	a=107471;b=537795;opcode=111;
			#100	a=988032;b=-355924;opcode=010;
			#100	a=5254;b=-525573;opcode=001;
			#100	a=369022;b=791055;opcode=111;
			#100	a=323602;b=-464376;opcode=110;
			#100	a=700205;b=14394;opcode=000;
			#100	a=-802679;b=-919308;opcode=111;
			#100	a=-658777;b=-694294;opcode=110;
			#100	a=-912386;b=-62632;opcode=100;
			#100	a=-317059;b=325642;opcode=001;
			#100	a=-401258;b=295791;opcode=001;
			#100	a=831463;b=-160781;opcode=010;
			#100	a=437323;b=-464744;opcode=100;
			#100	a=681023;b=-290123;opcode=111;
			#100	a=52252;b=806433;opcode=111;
			#100	a=643082;b=-225153;opcode=000;
			#100	a=-449920;b=-186788;opcode=100;
			#100	a=293109;b=-325139;opcode=100;
			#100	a=720397;b=-826217;opcode=001;
			#100	a=841644;b=994068;opcode=001;
			#100	a=-734707;b=-213148;opcode=111;
			#100	a=612378;b=225535;opcode=001;
			#100	a=740847;b=969750;opcode=111;
			#100	a=177564;b=-302997;opcode=000;
			#100	a=-395805;b=385988;opcode=000;
			#100	a=-25723;b=-473944;opcode=000;
			#100	a=411094;b=-593608;opcode=111;
			#100	a=-837336;b=692546;opcode=100;
			#100	a=-988371;b=-351990;opcode=111;
			#100	a=723211;b=285570;opcode=110;
			#100	a=-399413;b=-585309;opcode=111;
			#100	a=780770;b=441711;opcode=000;
			#100	a=31442;b=78932;opcode=111;
			#100	a=352485;b=-246560;opcode=001;
			#100	a=593404;b=-52943;opcode=110;
			#100	a=-391332;b=-356493;opcode=001;
			#100	a=3500;b=741459;opcode=010;
			#100	a=604558;b=247666;opcode=111;
			#100	a=447721;b=-874186;opcode=000;
			#100	a=-772553;b=691715;opcode=111;
			#100	a=809249;b=9586;opcode=010;
			#100	a=-932739;b=254794;opcode=110;
			#100	a=174989;b=450172;opcode=100;
			#100	a=-273291;b=823831;opcode=001;
			#100	a=486877;b=36576;opcode=001;
			#100	a=676384;b=459536;opcode=100;
			#100	a=526514;b=-142720;opcode=110;
			#100	a=729482;b=783671;opcode=000;
			#100	a=293108;b=110421;opcode=010;
			#100	a=539608;b=-594172;opcode=000;
			#100	a=-105397;b=-313924;opcode=100;
			#100	a=-205230;b=10160;opcode=111;
			#100	a=-88177;b=397649;opcode=010;
			#100	a=853203;b=-947233;opcode=010;
			#100	a=-641044;b=-884884;opcode=000;
			#100	a=-412542;b=137412;opcode=000;
			#100	a=624446;b=409042;opcode=010;
			#100	a=63108;b=713765;opcode=010;
			#100	a=-874925;b=-602870;opcode=000;
			#100	a=203091;b=-744664;opcode=111;
			#100	a=-919032;b=394598;opcode=100;
			#100	a=713031;b=-769175;opcode=100;
			#100	a=-833638;b=90622;opcode=000;
			#100	a=-576401;b=-555257;opcode=111;
			#100	a=724386;b=74998;opcode=001;
			#100	a=237221;b=-701464;opcode=110;
			#100	a=677679;b=95254;opcode=110;
			#100	a=-506494;b=116712;opcode=001;
			#100	a=90717;b=71571;opcode=010;
			#100	a=872970;b=-45100;opcode=100;
			#100	a=-33581;b=878368;opcode=100;
			#100	a=489152;b=639822;opcode=110;
			#100	a=943699;b=943454;opcode=110;
			#100	a=214107;b=577914;opcode=110;
			#100	a=369860;b=273981;opcode=110;
			#100	a=124445;b=-714524;opcode=001;
			#100	a=-988777;b=446229;opcode=001;
			#100	a=974832;b=803939;opcode=001;
			#100	a=-597343;b=-426717;opcode=001;
			#100	a=156858;b=-640176;opcode=100;
			#100	a=45153;b=-385776;opcode=010;
			#100	a=631255;b=959969;opcode=001;
			#100	a=-957025;b=212626;opcode=100;
			#100	a=665327;b=-820041;opcode=000;
			#100	a=188539;b=168627;opcode=110;
			#100	a=-182112;b=-710929;opcode=110;
			#100	a=-249095;b=870109;opcode=010;
			#100	a=831507;b=627601;opcode=110;
			#100	a=-127421;b=987885;opcode=001;
			#100	a=-665833;b=-920482;opcode=000;
			#100	a=913193;b=-562303;opcode=111;
			#100	a=-984488;b=-720780;opcode=111;
			#100	a=-859638;b=604792;opcode=110;
			#100	a=249130;b=-205541;opcode=010;
			#100	a=966209;b=-707483;opcode=100;
			#100	a=999040;b=-897321;opcode=010;
			#100	a=185252;b=-710730;opcode=000;
			#100	a=358873;b=-397916;opcode=000;
			#100	a=-195033;b=-435961;opcode=110;
			#100	a=-591599;b=569825;opcode=111;
			#100	a=202340;b=934050;opcode=010;
			#100	a=-198009;b=-30630;opcode=010;
			#100	a=-201947;b=22803;opcode=001;
			#100	a=571952;b=147699;opcode=010;
			#100	a=803084;b=-988727;opcode=110;
			#100	a=639691;b=-916249;opcode=001;
			#100	a=182851;b=290295;opcode=100;
			#100	a=719638;b=-11317;opcode=111;
			#100	a=-225554;b=-153364;opcode=100;
			#100	a=-727276;b=-958029;opcode=000;
			#100	a=399227;b=-721237;opcode=100;
			#100	a=341745;b=-841569;opcode=111;
			#100	a=148239;b=517378;opcode=110;
			#100	a=-426239;b=-313279;opcode=001;
			#100	a=671657;b=-547611;opcode=111;
			#100	a=-416001;b=-77852;opcode=010;
			#100	a=-738292;b=-980026;opcode=100;
			#100	a=-584940;b=-410526;opcode=100;
			#100	a=-379025;b=-328092;opcode=001;
			#100	a=-442024;b=-462468;opcode=000;
			#100	a=-888015;b=-364059;opcode=000;
			#100	a=212781;b=177062;opcode=100;
			#100	a=-166149;b=256814;opcode=100;
			#100	a=798674;b=-346130;opcode=000;
			#100	a=-610038;b=200649;opcode=100;
			#100	a=-147244;b=-131392;opcode=110;
			#100	a=-453085;b=-104838;opcode=100;
			#100	a=686223;b=-84930;opcode=111;
			#100	a=423971;b=-497266;opcode=001;
			#100	a=953178;b=68602;opcode=100;
			#100	a=-759120;b=208200;opcode=001;
			#100	a=-481575;b=-79110;opcode=010;
			#100	a=272034;b=561695;opcode=110;
			#100	a=599566;b=-317726;opcode=001;
			#100	a=-788328;b=-447580;opcode=000;
			#100	a=-249015;b=354477;opcode=001;
			#100	a=112118;b=-96856;opcode=000;
			#100	a=38834;b=544556;opcode=110;
			#100	a=974086;b=414326;opcode=001;
			#100	a=988946;b=-194809;opcode=001;
			#100	a=856222;b=712354;opcode=111;
			#100	a=805063;b=12774;opcode=010;
			#100	a=-513191;b=336478;opcode=100;
			#100	a=-229400;b=599356;opcode=100;
			#100	a=-421064;b=328421;opcode=001;
			#100	a=-988762;b=557166;opcode=110;
			#100	a=-403526;b=-224458;opcode=100;
			#100	a=834702;b=-801943;opcode=100;
			#100	a=279648;b=-295684;opcode=001;
			#100	a=-280773;b=-30687;opcode=111;
			#100	a=-883302;b=-625102;opcode=100;
			#100	a=355453;b=-799181;opcode=001;
			#100	a=661782;b=-839097;opcode=000;
			#100	a=-369144;b=-579381;opcode=010;
			#100	a=-696263;b=-771551;opcode=111;
			#100	a=205518;b=-967092;opcode=000;
			#100	a=844769;b=-125445;opcode=100;
			#100	a=226675;b=-261561;opcode=110;
			#100	a=629470;b=72688;opcode=001;
			#100	a=-47092;b=669034;opcode=001;
			#100	a=-475489;b=257903;opcode=110;
			#100	a=-670829;b=72803;opcode=111;
			#100	a=-305922;b=-731737;opcode=111;
			#100	a=60072;b=-574113;opcode=010;
			#100	a=-656860;b=582432;opcode=100;
			#100	a=-57149;b=-753586;opcode=111;
			#100	a=-37190;b=-229388;opcode=111;
			#100	a=242087;b=945463;opcode=000;
			#100	a=-499212;b=-231961;opcode=100;
			#100	a=335317;b=254798;opcode=100;
			#100	a=-545400;b=-935023;opcode=110;
			#100	a=-958706;b=809329;opcode=100;
			#100	a=-89057;b=-896626;opcode=111;
			#100	a=-282746;b=-482693;opcode=001;
			#100	a=312891;b=732481;opcode=001;
			#100	a=390203;b=-850964;opcode=100;
			#100	a=271563;b=-725579;opcode=100;
			#100	a=-152400;b=-775178;opcode=001;
			#100	a=-453508;b=420738;opcode=111;
			#100	a=72709;b=431728;opcode=100;
			#100	a=824199;b=479900;opcode=100;
			#100	a=503194;b=-203606;opcode=001;
			#100	a=-331584;b=-393201;opcode=010;
			#100	a=-560799;b=-925739;opcode=001;
			#100	a=694350;b=-577701;opcode=110;
			#100	a=130485;b=-24408;opcode=010;
			#100	a=-489021;b=-470027;opcode=111;
			#100	a=87002;b=245253;opcode=100;
			#100	a=-389087;b=-245362;opcode=010;
			#100	a=153715;b=489823;opcode=100;
			#100	a=186567;b=-606371;opcode=110;
			#100	a=141743;b=-786497;opcode=010;
			#100	a=123750;b=-931211;opcode=001;
			#100	a=-500125;b=-109823;opcode=001;
			#100	a=806433;b=-649797;opcode=100;
			#100	a=-897563;b=-430412;opcode=000;
			#100	a=623178;b=-896982;opcode=001;
			#100	a=-725190;b=858037;opcode=111;
			#100	a=-412842;b=-793526;opcode=000;
			#100	a=-912352;b=577821;opcode=000;
			#100	a=515379;b=-769502;opcode=010;
			#100	a=-500075;b=-255305;opcode=110;
			#100	a=516506;b=-23685;opcode=001;
			#100	a=-479275;b=983354;opcode=100;
			#100	a=285942;b=-304649;opcode=111;
			#100	a=671817;b=-621675;opcode=010;
			#100	a=-141989;b=-32949;opcode=100;
			#100	a=910727;b=-6636;opcode=000;
			#100	a=568156;b=-200547;opcode=001;
			#100	a=-638366;b=-426554;opcode=001;
			#100	a=191156;b=582353;opcode=100;
			#100	a=738527;b=812139;opcode=000;
			#100	a=653176;b=-518465;opcode=100;
			#100	a=-790678;b=-811033;opcode=001;
			#100	a=618107;b=-521224;opcode=100;
			#100	a=794248;b=-437806;opcode=010;
			#100	a=296234;b=950961;opcode=010;
			#100	a=-764424;b=-254933;opcode=010;
			#100	a=-591197;b=-734104;opcode=000;
			#100	a=652900;b=-106840;opcode=010;
			#100	a=54395;b=811249;opcode=001;
			#100	a=279043;b=152256;opcode=110;
			#100	a=-255587;b=533709;opcode=111;
			#100	a=766183;b=-280701;opcode=000;
			#100	a=563414;b=99599;opcode=010;
			#100	a=-163550;b=568310;opcode=111;
			#100	a=945935;b=624028;opcode=111;
			#100	a=262439;b=828912;opcode=100;
			#100	a=-141631;b=603533;opcode=001;
			#100	a=384680;b=-791708;opcode=111;
			#100	a=-577547;b=-264301;opcode=001;
			#100	a=764256;b=356339;opcode=010;
			#100	a=116596;b=-914831;opcode=100;
			#100	a=583043;b=430606;opcode=111;
			#100	a=343367;b=243042;opcode=100;
			#100	a=981022;b=-516438;opcode=000;
			#100	a=-284523;b=816408;opcode=001;
			#100	a=948567;b=-721684;opcode=111;
			#100	a=147648;b=972645;opcode=110;
			#100	a=-602040;b=110743;opcode=010;
			#100	a=-220765;b=-149144;opcode=110;
			#100	a=-888001;b=-689258;opcode=000;
			#100	a=706368;b=117964;opcode=100;
			#100	a=-752638;b=-377476;opcode=010;
			#100	a=47163;b=662062;opcode=001;
			#100	a=-237560;b=804628;opcode=111;
			#100	a=-857270;b=-797898;opcode=111;
			#100	a=-12416;b=94214;opcode=010;
			#100	a=-267758;b=-363054;opcode=000;
			#100	a=786175;b=180442;opcode=100;
			#100	a=-102370;b=-428253;opcode=111;
			#100	a=-198754;b=856782;opcode=001;
			#100	a=932036;b=755641;opcode=100;
			#100	a=-820820;b=-440953;opcode=001;
			#100	a=939319;b=586002;opcode=100;
			#100	a=405021;b=194804;opcode=111;
			#100	a=-54227;b=-500024;opcode=111;
			#100	a=-253082;b=-362725;opcode=100;
			#100	a=-979676;b=32227;opcode=100;
			#100	a=-773053;b=104797;opcode=000;
			#100	a=867478;b=-209780;opcode=111;
			#100	a=-814599;b=-284877;opcode=001;
			#100	a=341929;b=3705;opcode=000;
			#100	a=594119;b=726774;opcode=010;
			#100	a=306771;b=-627963;opcode=111;
			#100	a=146598;b=-78348;opcode=001;
			#100	a=-373322;b=-22569;opcode=110;
			#100	a=-635538;b=960713;opcode=110;
			#100	a=-876325;b=-943611;opcode=000;
			#100	a=979563;b=707746;opcode=001;
			#100	a=-625481;b=506990;opcode=000;
			#100	a=795348;b=407995;opcode=000;
			#100	a=-414045;b=853992;opcode=000;
			#100	a=112470;b=461816;opcode=000;
			#100	a=780143;b=-835367;opcode=000;
			#100	a=212532;b=-644618;opcode=001;
			#100	a=-458085;b=9522;opcode=000;
			#100	a=687966;b=169406;opcode=000;
			#100	a=-714098;b=-425641;opcode=010;
			#100	a=50941;b=394719;opcode=010;
			#100	a=111129;b=-350871;opcode=100;
			#100	a=924242;b=-810861;opcode=010;
			#100	a=-721406;b=-587656;opcode=111;
			#100	a=-810807;b=393931;opcode=000;
			#100	a=-500302;b=297895;opcode=000;
			#100	a=723183;b=101413;opcode=100;
			#100	a=-127778;b=-746008;opcode=001;
			#100	a=-459544;b=17920;opcode=001;
			#100	a=864415;b=-773122;opcode=110;
			#100	a=263395;b=487877;opcode=010;
			#100	a=741604;b=-117930;opcode=001;
			#100	a=547390;b=-6398;opcode=111;
			#100	a=529647;b=547093;opcode=010;
			#100	a=-516381;b=-200335;opcode=111;
			#100	a=878829;b=-113239;opcode=111;
			#100	a=262448;b=493385;opcode=010;
			#100	a=-229342;b=754945;opcode=010;
			#100	a=535694;b=-604955;opcode=100;
			#100	a=349450;b=-719122;opcode=010;
			#100	a=265417;b=370283;opcode=100;
			#100	a=-80064;b=269677;opcode=110;
			#100	a=-460347;b=-589033;opcode=010;
			#100	a=-225469;b=-929338;opcode=010;
			#100	a=-828688;b=-617178;opcode=110;
			#100	a=717405;b=-753946;opcode=100;
			#100	a=-606499;b=452321;opcode=001;
			#100	a=-471943;b=251211;opcode=100;
			#100	a=-427235;b=-976254;opcode=000;
			#100	a=422082;b=-419917;opcode=001;
			#100	a=-777522;b=-84897;opcode=100;
			#100	a=-310884;b=-726931;opcode=110;
			#100	a=275339;b=-514352;opcode=010;
			#100	a=773951;b=-29348;opcode=001;
			#100	a=-45603;b=-547119;opcode=110;
			#100	a=-406110;b=29406;opcode=000;
			#100	a=-370921;b=-444134;opcode=010;
			#100	a=-134143;b=956824;opcode=000;
			#100	a=-137749;b=48817;opcode=010;
			#100	a=843996;b=979060;opcode=111;
			#100	a=-345211;b=828842;opcode=110;
			#100	a=981746;b=472270;opcode=001;
			#100	a=-575474;b=-6249;opcode=010;
			#100	a=602775;b=-20028;opcode=001;
			#100	a=-589586;b=89625;opcode=111;
			#100	a=367726;b=-232942;opcode=001;
			#100	a=-50357;b=-884139;opcode=110;
			#100	a=882406;b=-228700;opcode=000;
			#100	a=-30819;b=-642339;opcode=010;
			#100	a=-420758;b=-871385;opcode=100;
			#100	a=-555767;b=911357;opcode=110;
			#100	a=266782;b=866243;opcode=110;
			#100	a=876513;b=782265;opcode=001;
			#100	a=305997;b=355058;opcode=001;
			#100	a=249678;b=-673849;opcode=001;
			#100	a=-706151;b=308314;opcode=000;
			#100	a=490845;b=-461398;opcode=110;
			#100	a=123578;b=220929;opcode=100;
			#100	a=-125608;b=-355635;opcode=111;
			#100	a=574560;b=911490;opcode=000;
			#100	a=666360;b=-783353;opcode=010;
			#100	a=-42326;b=312622;opcode=000;
			#100	a=-433464;b=792053;opcode=100;
			#100	a=792126;b=-670575;opcode=100;
			#100	a=-812100;b=496924;opcode=010;
			#100	a=639096;b=-206529;opcode=010;
			#100	a=455862;b=399790;opcode=111;
			#100	a=-226920;b=637257;opcode=010;
			#100	a=395532;b=20693;opcode=001;
			#100	a=-216256;b=99721;opcode=001;
			#100	a=-261040;b=518542;opcode=110;
			#100	a=-298019;b=-787816;opcode=110;
			#100	a=50101;b=-261293;opcode=001;
			#100	a=577856;b=-672089;opcode=111;
			#100	a=-360909;b=-226144;opcode=111;
			#100	a=111229;b=-131068;opcode=001;
			#100	a=541065;b=-706862;opcode=001;
			#100	a=474855;b=779765;opcode=000;
			#100	a=-762491;b=675230;opcode=100;
			#100	a=-586324;b=-717919;opcode=001;
			#100	a=566323;b=35546;opcode=110;
			#100	a=-413376;b=603643;opcode=010;
			#100	a=-624281;b=-938338;opcode=110;
			#100	a=-110262;b=358115;opcode=100;
			#100	a=-619131;b=-241570;opcode=010;
			#100	a=-278471;b=372180;opcode=000;
			#100	a=714450;b=577325;opcode=010;
			#100	a=-150422;b=-801041;opcode=001;
			#100	a=772012;b=-304988;opcode=100;
			#100	a=-960160;b=-953874;opcode=001;
			#100	a=-408713;b=784360;opcode=100;
			#100	a=-476603;b=430237;opcode=100;
			#100	a=160510;b=-246648;opcode=111;
			#100	a=-196017;b=315951;opcode=111;
			#100	a=-703441;b=-654970;opcode=110;
			#100	a=-22925;b=-602366;opcode=010;
			#100	a=499613;b=-905175;opcode=001;
			#100	a=-945367;b=867932;opcode=111;
			#100	a=-689956;b=500820;opcode=001;
			#100	a=-329166;b=40638;opcode=010;
			#100	a=-136642;b=384477;opcode=010;
			#100	a=-986965;b=607605;opcode=100;
			#100	a=-384618;b=964163;opcode=001;
			#100	a=87801;b=468626;opcode=010;
			#100	a=-630295;b=357519;opcode=111;
			#100	a=-122636;b=-63112;opcode=110;
			#100	a=781573;b=-318090;opcode=010;
			#100	a=336888;b=92104;opcode=111;
			#100	a=958934;b=-76346;opcode=010;
			#100	a=580144;b=168841;opcode=111;
			#100	a=453199;b=671456;opcode=000;
			#100	a=611241;b=-245346;opcode=110;
			#100	a=-69276;b=-238355;opcode=111;
			#100	a=-127686;b=-902054;opcode=001;
			#100	a=-427894;b=79806;opcode=000;
			#100	a=179948;b=182231;opcode=001;
			#100	a=-981953;b=-84248;opcode=001;
			#100	a=921627;b=936657;opcode=100;
			#100	a=-268503;b=567801;opcode=100;
			#100	a=-361865;b=-866320;opcode=100;
			#100	a=136194;b=-472903;opcode=000;
			#100	a=-369670;b=-115095;opcode=010;
			#100	a=-401198;b=-251510;opcode=100;
			#100	a=-596437;b=612228;opcode=100;
			#100	a=-264213;b=633737;opcode=110;
			#100	a=587074;b=-134816;opcode=111;
			#100	a=748318;b=435921;opcode=010;
			#100	a=914578;b=-932777;opcode=010;
			#100	a=108012;b=151901;opcode=100;
			#100	a=-265731;b=821324;opcode=100;
			#100	a=711523;b=372805;opcode=100;
			#100	a=702069;b=755823;opcode=110;
			#100	a=-762853;b=760035;opcode=111;
			#100	a=-7355;b=-898395;opcode=001;
			#100	a=-691897;b=-850815;opcode=001;
			#100	a=-791564;b=-187485;opcode=111;
			#100	a=898087;b=619050;opcode=110;
			#100	a=-469528;b=-528256;opcode=110;
			#100	a=-208578;b=-431332;opcode=111;
			#100	a=265329;b=-288085;opcode=000;
			#100	a=777091;b=616657;opcode=000;
			#100	a=316314;b=-839313;opcode=000;
			#100	a=553889;b=-193363;opcode=010;
			#100	a=-341416;b=-58350;opcode=001;
			#100	a=-726256;b=-251086;opcode=100;
			#100	a=-914198;b=-904985;opcode=001;
			#100	a=128472;b=595688;opcode=000;
			#100	a=-676007;b=-72509;opcode=000;
			#100	a=-952692;b=320329;opcode=001;
			#100	a=-872092;b=671343;opcode=010;
			#100	a=791130;b=-75149;opcode=001;
			#100	a=-480352;b=333060;opcode=110;
			#100	a=-573968;b=452977;opcode=111;
			#100	a=-214742;b=828601;opcode=000;
			#100	a=-431952;b=-902333;opcode=111;
			#100	a=295831;b=-180631;opcode=111;
			#100	a=-22291;b=551186;opcode=111;
			#100	a=571740;b=-772571;opcode=100;
			#100	a=7320;b=-681224;opcode=111;
			#100	a=-444083;b=509821;opcode=001;
			#100	a=-588657;b=-802988;opcode=100;
			#100	a=-973739;b=-290438;opcode=111;
			#100	a=-838772;b=-476980;opcode=111;
			#100	a=-935878;b=668054;opcode=010;
			#100	a=125938;b=-827446;opcode=010;
			#100	a=-668720;b=-509430;opcode=001;
			#100	a=563905;b=153642;opcode=110;
			#100	a=392032;b=-466985;opcode=000;
			#100	a=39415;b=997192;opcode=000;
			#100	a=-229712;b=789117;opcode=001;
			#100	a=256129;b=-765781;opcode=111;
			#100	a=-810719;b=-472078;opcode=010;
			#100	a=966212;b=-533141;opcode=100;
			#100	a=-174252;b=-654469;opcode=000;
			#100	a=216763;b=186883;opcode=010;
			#100	a=-431196;b=-794468;opcode=001;
			#100	a=-699458;b=-470948;opcode=010;
			#100	a=-114474;b=558332;opcode=000;
			#100	a=8410;b=-711219;opcode=001;
			#100	a=-629166;b=-196070;opcode=000;
			#100	a=-393714;b=620465;opcode=001;
			#100	a=-737699;b=508527;opcode=111;
			#100	a=-368686;b=-681473;opcode=110;
			#100	a=237617;b=-881831;opcode=010;
			#100	a=-326217;b=911679;opcode=100;
			#100	a=-206958;b=554734;opcode=110;
			#100	a=-480693;b=514329;opcode=010;
			#100	a=-109397;b=143098;opcode=010;
			#100	a=103941;b=165868;opcode=000;
			#100	a=870789;b=60133;opcode=010;
			#100	a=-621966;b=-763593;opcode=000;
			#100	a=834406;b=800346;opcode=010;
			#100	a=764517;b=-214067;opcode=111;
			#100	a=616533;b=-406619;opcode=100;
			#100	a=-557841;b=-218455;opcode=110;
			#100	a=-809649;b=-413716;opcode=001;
			#100	a=-361915;b=804845;opcode=111;
			#100	a=257007;b=787757;opcode=110;
			#100	a=-811346;b=-113484;opcode=111;
			#100	a=-22940;b=-933621;opcode=010;
			#100	a=-342357;b=-397874;opcode=000;
			#100	a=-851006;b=707651;opcode=001;
			#100	a=-354003;b=-532855;opcode=001;
			#100	a=682663;b=-303946;opcode=111;
			#100	a=-465677;b=-220363;opcode=010;
			#100	a=846830;b=866854;opcode=001;
			#100	a=158494;b=-225719;opcode=000;
			#100	a=-363738;b=149226;opcode=001;
			#100	a=476809;b=136440;opcode=111;
			#100	a=-455285;b=-73912;opcode=001;
			#100	a=-344082;b=-104715;opcode=001;
			#100	a=899658;b=-378317;opcode=000;
			#100	a=-206218;b=519468;opcode=010;
			#100	a=934613;b=-131350;opcode=110;
			#100	a=-518499;b=-671293;opcode=001;
			#100	a=645569;b=-227837;opcode=111;
			#100	a=-374182;b=-283725;opcode=010;
			#100	a=729663;b=566580;opcode=111;
			#100	a=714819;b=-142375;opcode=001;
			#100	a=-200880;b=807424;opcode=010;
			#100	a=504403;b=-389518;opcode=000;
			#100	a=-491632;b=370650;opcode=111;
			#100	a=448389;b=-852152;opcode=001;
			#100	a=256162;b=-791501;opcode=000;
			#100	a=-676224;b=719548;opcode=111;
			#100	a=-253817;b=-818427;opcode=010;
			#100	a=-744625;b=499909;opcode=111;
			#100	a=-283511;b=-479859;opcode=111;
			#100	a=-127555;b=932143;opcode=110;
			#100	a=390867;b=-241840;opcode=110;
			#100	a=413246;b=-35364;opcode=110;
			#100	a=-326476;b=-246377;opcode=111;
			#100	a=120157;b=519757;opcode=100;
			#100	a=265690;b=385894;opcode=001;
			#100	a=157635;b=-166303;opcode=110;
			#100	a=250897;b=-72777;opcode=010;
			#100	a=-612941;b=-340307;opcode=100;
			#100	a=-977341;b=756626;opcode=110;
			#100	a=852171;b=-161762;opcode=010;
			#100	a=-86958;b=-791118;opcode=100;
			#100	a=118889;b=592283;opcode=001;
			#100	a=110137;b=146177;opcode=010;
			#100	a=618164;b=-108153;opcode=010;
			#100	a=-895481;b=-694982;opcode=110;
			#100	a=827309;b=336159;opcode=001;
			#100	a=846690;b=260985;opcode=001;
			#100	a=216596;b=97675;opcode=111;
			#100	a=238210;b=982386;opcode=001;
			#100	a=-448193;b=942956;opcode=000;
			#100	a=902949;b=802754;opcode=010;
			#100	a=-808123;b=-923817;opcode=100;
			#100	a=842551;b=134470;opcode=111;
			#100	a=309432;b=-106096;opcode=100;
			#100	a=-407397;b=548303;opcode=110;
			#100	a=158931;b=-912794;opcode=000;
			#100	a=-671842;b=23823;opcode=001;
			#100	a=872730;b=435244;opcode=010;
			#100	a=587201;b=204617;opcode=000;
			#100	a=-301192;b=505936;opcode=111;
			#100	a=-549037;b=-344471;opcode=111;
			#100	a=-174902;b=-145740;opcode=111;
			#100	a=163039;b=742546;opcode=110;
			#100	a=-543367;b=-698508;opcode=110;
			#100	a=-242034;b=747229;opcode=111;
			#100	a=-293736;b=976125;opcode=111;
			#100	a=970015;b=12704;opcode=110;
			#100	a=524987;b=573891;opcode=001;
			#100	a=-482063;b=-320024;opcode=110;
			#100	a=-608448;b=744987;opcode=100;
			#100	a=840022;b=-749648;opcode=111;
			#100	a=984513;b=529456;opcode=110;
			#100	a=31626;b=452460;opcode=111;
			#100	a=536779;b=-159663;opcode=000;
			#100	a=-536413;b=-843;opcode=010;
			#100	a=-216324;b=-803633;opcode=111;
			#100	a=-647866;b=-884250;opcode=000;
			#100	a=164195;b=-748199;opcode=100;
			#100	a=-222295;b=497316;opcode=001;
			#100	a=827161;b=903896;opcode=000;
			#100	a=-735232;b=10990;opcode=001;
			#100	a=595236;b=-335979;opcode=100;
			#100	a=-700389;b=-183783;opcode=001;
			#100	a=301152;b=978520;opcode=100;
			#100	a=-511997;b=-646052;opcode=111;
			#100	a=287362;b=321347;opcode=001;
			#100	a=-803556;b=286158;opcode=111;
			#100	a=263408;b=953732;opcode=001;
			#100	a=961333;b=90486;opcode=111;
			#100	a=217971;b=-675064;opcode=111;
			#100	a=-618592;b=-159052;opcode=000;
			#100	a=393922;b=-812623;opcode=001;
			#100	a=386017;b=265096;opcode=010;
			#100	a=-875049;b=940749;opcode=000;
			#100	a=302196;b=589788;opcode=100;
			#100	a=-248311;b=-592535;opcode=100;
			#100	a=-512482;b=339015;opcode=111;
			#100	a=354504;b=-675024;opcode=001;
			#100	a=255026;b=338437;opcode=000;
			#100	a=-384444;b=-217023;opcode=010;
			#100	a=281155;b=-120710;opcode=110;
			#100	a=-998071;b=428143;opcode=000;
			#100	a=-444923;b=-282720;opcode=100;
			#100	a=289884;b=-568482;opcode=001;
			#100	a=-890114;b=561195;opcode=111;
			#100	a=-278076;b=-47234;opcode=010;
			#100	a=212038;b=515769;opcode=001;
			#100	a=462447;b=193456;opcode=010;
			#100	a=-171547;b=-139078;opcode=111;
			#100	a=303552;b=225770;opcode=111;
			#100	a=762890;b=-920764;opcode=000;
			#100	a=-104533;b=92151;opcode=111;
			#100	a=262674;b=637734;opcode=010;
			#100	a=951681;b=109715;opcode=100;
			#100	a=326716;b=-262585;opcode=100;
			#100	a=166548;b=657572;opcode=110;
			#100	a=-135073;b=262471;opcode=001;
			#100	a=670071;b=849805;opcode=111;
			#100	a=460239;b=-835152;opcode=000;
			#100	a=613835;b=-121280;opcode=100;
			#100	a=-273983;b=-665565;opcode=110;
			#100	a=-57661;b=-180403;opcode=000;
			#100	a=-960697;b=-44410;opcode=110;
			#100	a=62859;b=357838;opcode=110;
			#100	a=908295;b=-717534;opcode=111;
			#100	a=-666680;b=622876;opcode=111;
			#100	a=-259672;b=-456293;opcode=110;
			#100	a=452378;b=185420;opcode=001;
			#100	a=-893457;b=-717755;opcode=110;
			#100	a=581640;b=-89519;opcode=001;
			#100	a=764379;b=9561;opcode=010;
			#100	a=-509570;b=-842183;opcode=010;
			#100	a=-662117;b=505462;opcode=100;
			#100	a=-692392;b=-851059;opcode=100;
			#100	a=111340;b=-941402;opcode=001;
			#100	a=101914;b=940282;opcode=010;
			#100	a=-36191;b=191710;opcode=111;
			#100	a=-102210;b=952152;opcode=100;
			#100	a=-438098;b=476067;opcode=001;
			#100	a=-656311;b=64368;opcode=111;
			#100	a=-540371;b=786385;opcode=111;
			#100	a=-577570;b=420620;opcode=001;
			#100	a=269882;b=-814149;opcode=110;
			#100	a=-783230;b=-695896;opcode=001;
			#100	a=-745443;b=376689;opcode=001;
			#100	a=280435;b=992859;opcode=001;
			#100	a=-25070;b=-406024;opcode=111;
			#100	a=-925207;b=-556771;opcode=100;
			#100	a=-593917;b=838390;opcode=000;
			#100	a=-967620;b=412268;opcode=110;
			#100	a=-187632;b=780301;opcode=110;
			#100	a=720270;b=-588133;opcode=111;
			#100	a=-736540;b=140047;opcode=110;
			#100	a=-58325;b=-601285;opcode=111;
			#100	a=170822;b=388702;opcode=110;
			#100	a=710185;b=-625753;opcode=000;
			#100	a=-788762;b=-519380;opcode=001;
			#100	a=-852233;b=639569;opcode=000;
			#100	a=943108;b=839502;opcode=111;
			#100	a=-623658;b=-324177;opcode=010;
			#100	a=-722183;b=-495232;opcode=010;
			#100	a=-25441;b=-294616;opcode=010;
			#100	a=325451;b=398243;opcode=100;
			#100	a=-945899;b=-428019;opcode=111;
			#100	a=425722;b=-258207;opcode=001;
			#100	a=228262;b=432442;opcode=100;
			#100	a=940906;b=-842416;opcode=001;
			#100	a=-555832;b=633783;opcode=100;
			#100	a=218644;b=418384;opcode=010;
			#100	a=-221895;b=369574;opcode=010;
			#100	a=-235262;b=-483019;opcode=001;
			#100	a=406377;b=5937;opcode=110;
			#100	a=186475;b=-478278;opcode=100;
			#100	a=81648;b=-372783;opcode=100;
			#100	a=984740;b=-453665;opcode=000;
			#100	a=-174334;b=-439851;opcode=010;
			#100	a=-800935;b=74383;opcode=010;
			#100	a=-243502;b=-692731;opcode=100;
			#100	a=-308696;b=-968588;opcode=001;
			#100	a=-327526;b=-563342;opcode=111;
			#100	a=733756;b=-471216;opcode=100;
			#100	a=628613;b=664495;opcode=111;
			#100	a=187840;b=511560;opcode=110;
			#100	a=506770;b=4629;opcode=100;
			#100	a=325126;b=-563445;opcode=010;
			#100	a=547370;b=15993;opcode=111;
			#100	a=23149;b=463084;opcode=111;
			#100	a=-472261;b=-5095;opcode=010;
			#100	a=251625;b=871541;opcode=010;
			#100	a=-165932;b=642341;opcode=010;
			#100	a=-558260;b=386577;opcode=001;
			#100	a=-59171;b=871552;opcode=000;
			#100	a=772398;b=-450971;opcode=000;
			#100	a=-127354;b=-682422;opcode=110;
			#100	a=-400178;b=447602;opcode=001;
			#100	a=-667831;b=-288751;opcode=010;
			#100	a=368580;b=-533986;opcode=001;
			#100	a=-974829;b=-857814;opcode=111;
			#100	a=630208;b=846497;opcode=111;
			#100	a=-129677;b=-721285;opcode=100;
			#100	a=-209065;b=276049;opcode=010;
			#100	a=-376526;b=-970051;opcode=100;
			#100	a=241360;b=-643185;opcode=100;
			#100	a=839605;b=518391;opcode=110;
			#100	a=-348242;b=433650;opcode=110;
			#100	a=-325489;b=707141;opcode=100;
			#100	a=-55935;b=939299;opcode=000;
			#100	a=-614143;b=134839;opcode=001;
			#100	a=-340176;b=-230840;opcode=010;
			#100	a=-156782;b=456506;opcode=110;
			#100	a=957794;b=968759;opcode=110;
			#100	a=-403922;b=-554801;opcode=010;
			#100	a=63696;b=-839375;opcode=111;
			#100	a=-980413;b=886515;opcode=110;
			#100	a=320056;b=227301;opcode=100;
			#100	a=-645487;b=-45848;opcode=001;
			#100	a=422139;b=-546292;opcode=000;
			#100	a=927353;b=973097;opcode=111;
			#100	a=521310;b=-965000;opcode=010;
			#100	a=350849;b=-827155;opcode=010;
			#100	a=-225633;b=-257618;opcode=111;
			#100	a=254950;b=-412443;opcode=000;
			#100	a=318035;b=-145965;opcode=100;
			#100	a=506694;b=-965173;opcode=100;
			#100	a=-472723;b=-583251;opcode=001;
			#100	a=327889;b=-130441;opcode=111;
			#100	a=-620876;b=134671;opcode=111;
			#100	a=-428209;b=-154946;opcode=001;
			#100	a=28302;b=242529;opcode=000;
			#100	a=212667;b=225767;opcode=100;
			#100	a=-326176;b=-780456;opcode=010;
			#100	a=664684;b=-520091;opcode=110;
			#100	a=-641527;b=-497087;opcode=110;
			#100	a=-274163;b=-375291;opcode=010;
			#100	a=-778405;b=180290;opcode=010;
			#100	a=762551;b=-802464;opcode=110;
			#100	a=225650;b=-102369;opcode=110;
			#100	a=-750420;b=781958;opcode=110;
			#100	a=-742866;b=-778839;opcode=000;
			#100	a=610796;b=-604524;opcode=111;
			#100	a=320794;b=-530805;opcode=100;
			#100	a=621486;b=771131;opcode=100;
			#100	a=-241507;b=936832;opcode=010;
			#100	a=481351;b=845282;opcode=001;
			#100	a=263334;b=-462496;opcode=100;
			#100	a=-886616;b=480052;opcode=100;
			#100	a=-445543;b=83140;opcode=010;
			#100	a=591171;b=-539825;opcode=010;
			#100	a=650688;b=-433593;opcode=111;
			#100	a=861891;b=-165904;opcode=000;
			#100	a=-586801;b=-8761;opcode=000;
			#100	a=744752;b=453967;opcode=111;
			#100	a=658538;b=618172;opcode=000;
			#100	a=-879280;b=509204;opcode=001;
			#100	a=307175;b=163974;opcode=111;
			#100	a=-167076;b=156951;opcode=110;
			#100	a=54488;b=-370847;opcode=110;
			#100	a=910744;b=105541;opcode=100;
			#100	a=-652778;b=346655;opcode=111;
			#100	a=76604;b=841766;opcode=000;
			#100	a=575818;b=-861801;opcode=110;
			#100	a=871554;b=-450106;opcode=001;
			#100	a=668562;b=-379877;opcode=111;
			#100	a=-696863;b=587266;opcode=110;
			#100	a=-911868;b=493381;opcode=110;
			#100	a=-431028;b=128218;opcode=111;
			#100	a=660825;b=-793946;opcode=010;
			#100	a=227017;b=-636677;opcode=100;
			#100	a=-745849;b=475871;opcode=110;
			#100	a=-784564;b=412823;opcode=100;
			#100	a=881567;b=-987313;opcode=010;
			#100	a=-871767;b=245816;opcode=010;
			#100	a=-941787;b=-308844;opcode=000;
			#100	a=242985;b=-275122;opcode=000;
			#100	a=-104197;b=-979730;opcode=110;
			#100	a=182734;b=-979234;opcode=010;
			#100	a=-95118;b=235527;opcode=010;
			#100	a=-452177;b=-188801;opcode=000;
			#100	a=-321288;b=-126783;opcode=000;
			#100	a=-317648;b=-803308;opcode=111;
			#100	a=-437158;b=-821353;opcode=000;
			#100	a=875169;b=811175;opcode=001;
			#100	a=263571;b=-794862;opcode=100;
			#100	a=-45313;b=-887024;opcode=110;
			#100	a=415980;b=-450759;opcode=111;
			#100	a=9941;b=461339;opcode=001;
			#100	a=392770;b=-52245;opcode=111;
			#100	a=813647;b=331396;opcode=110;
			#100	a=-349465;b=-389932;opcode=010;
			#100	a=-561241;b=-779107;opcode=001;
			#100	a=-361566;b=605478;opcode=001;
			#100	a=-894038;b=282729;opcode=010;
			#100	a=-611403;b=310530;opcode=001;
			#100	a=93516;b=-27848;opcode=111;
			#100	a=-130179;b=-918741;opcode=010;
			#100	a=-745114;b=172319;opcode=000;
			#100	a=146044;b=-211669;opcode=000;
			#100	a=1740;b=641518;opcode=001;
			#100	a=448368;b=653801;opcode=110;
			#100	a=-195410;b=-827577;opcode=111;
			#100	a=-772752;b=410773;opcode=010;
			#100	a=864769;b=-763517;opcode=010;
			#100	a=958454;b=268650;opcode=000;
			#100	a=-888966;b=-628604;opcode=110;
			#100	a=-911137;b=-29454;opcode=000;
			#100	a=696099;b=-53643;opcode=111;
			#100	a=-759622;b=-415020;opcode=111;
			#100	a=679791;b=372019;opcode=001;
			#100	a=473449;b=-885596;opcode=110;
			#100	a=-238406;b=-902186;opcode=001;
			#100	a=667927;b=97970;opcode=010;
			#100	a=972524;b=-273782;opcode=001;
			#100	a=-866805;b=-789195;opcode=100;
			#100	a=158239;b=-463485;opcode=000;
			#100	a=1610;b=361039;opcode=010;
			#100	a=-776981;b=549029;opcode=001;
			#100	a=800883;b=206535;opcode=000;
			#100	a=110708;b=-438618;opcode=100;
			#100	a=842710;b=-126813;opcode=010;
			#100	a=-408357;b=-165398;opcode=111;
			#100	a=-625184;b=-334654;opcode=100;
			#100	a=679741;b=-313493;opcode=111;
			#100	a=404043;b=182232;opcode=010;
			#100	a=51321;b=128533;opcode=010;
			#100	a=383212;b=-11589;opcode=111;
			#100	a=-939287;b=490199;opcode=100;
			#100	a=-547789;b=597285;opcode=111;
			#100	a=-455155;b=-206219;opcode=001;
			#100	a=-452649;b=-945831;opcode=000;
			#100	a=-267371;b=-337803;opcode=000;
			#100	a=858038;b=480767;opcode=111;
			#100	a=-765857;b=-534373;opcode=110;
			#100	a=-416690;b=141610;opcode=001;
			#100	a=746160;b=-35895;opcode=000;
			#100	a=-139037;b=-183517;opcode=111;
			#100	a=695043;b=-96296;opcode=001;
			#100	a=763985;b=-412522;opcode=001;
			#100	a=-245400;b=451142;opcode=111;
			#100	a=-107761;b=289224;opcode=110;
			#100	a=972764;b=-490224;opcode=100;
			#100	a=-514504;b=636569;opcode=110;
			#100	a=-877039;b=-290587;opcode=000;
			#100	a=449174;b=-44000;opcode=111;
			#100	a=-263825;b=-661999;opcode=111;
			#100	a=876501;b=680964;opcode=010;
			#100	a=985027;b=-648318;opcode=110;
			#100	a=864157;b=-417363;opcode=010;
			#100	a=438374;b=628835;opcode=000;
			#100	a=31102;b=460605;opcode=111;
			#100	a=-366046;b=-669152;opcode=100;
			#100	a=-648162;b=-308116;opcode=110;
			#100	a=-639433;b=-510661;opcode=110;
			#100	a=-588511;b=-732941;opcode=000;
			#100	a=910637;b=-135523;opcode=000;
			#100	a=341306;b=-446196;opcode=100;
			#100	a=709731;b=613158;opcode=110;
			#100	a=-654720;b=-742062;opcode=111;
			#100	a=369929;b=-416117;opcode=010;
			#100	a=675903;b=700012;opcode=010;
			#100	a=472745;b=241418;opcode=001;
			#100	a=-966408;b=27459;opcode=110;
			#100	a=-64954;b=778536;opcode=001;
			#100	a=147221;b=-180881;opcode=100;
			#100	a=-578835;b=-235317;opcode=110;
			#100	a=289585;b=-502285;opcode=000;
			#100	a=120408;b=271473;opcode=110;
			#100	a=-6011;b=-449483;opcode=000;
			#100	a=538595;b=-148223;opcode=010;
			#100	a=402135;b=316120;opcode=110;
			#100	a=167963;b=967840;opcode=111;
			#100	a=185714;b=392588;opcode=000;
			#100	a=89477;b=-696325;opcode=010;
			#100	a=960906;b=-465792;opcode=100;
			#100	a=435967;b=788589;opcode=010;
			#100	a=538169;b=998731;opcode=100;
			#100	a=-36070;b=-808634;opcode=110;
			#100	a=46976;b=-914149;opcode=100;
			#100	a=-196866;b=-295733;opcode=010;
			#100	a=-243874;b=323841;opcode=110;
			#100	a=902104;b=-839087;opcode=100;
			#100	a=-659292;b=-420167;opcode=000;
			#100	a=-445640;b=-120861;opcode=100;
			#100	a=664027;b=-140101;opcode=110;
			#100	a=520795;b=283167;opcode=010;
			#100	a=-156240;b=336051;opcode=100;
			#100	a=514769;b=-12694;opcode=110;
			#100	a=93179;b=-891515;opcode=000;
			#100	a=-749391;b=149815;opcode=100;
			#100	a=-547130;b=-953800;opcode=010;
			#100	a=78757;b=594581;opcode=010;
			#100	a=-457808;b=-962464;opcode=000;
			#100	a=393780;b=136797;opcode=110;
			#100	a=-105203;b=651024;opcode=001;
			#100	a=621270;b=323616;opcode=001;
			#100	a=772665;b=12095;opcode=001;
			#100	a=476021;b=837827;opcode=111;
			#100	a=-573374;b=-839118;opcode=001;
			#100	a=251552;b=347337;opcode=010;
			#100	a=6916;b=813905;opcode=100;
			#100	a=-705735;b=-165073;opcode=111;
			#100	a=438675;b=353996;opcode=010;
			#100	a=158998;b=165953;opcode=110;
			#100	a=62654;b=539431;opcode=000;
			#100	a=256684;b=-677099;opcode=010;
			#100	a=-459038;b=773882;opcode=001;
			#100	a=-893984;b=791172;opcode=100;
			#100	a=75945;b=-252652;opcode=100;
			#100	a=-663595;b=598380;opcode=111;
			#100	a=211073;b=-945336;opcode=000;
			#100	a=-850914;b=-289498;opcode=010;
			#100	a=-332786;b=-345564;opcode=110;
			#100	a=-465602;b=783957;opcode=110;
			#100	a=834174;b=-553240;opcode=100;
			#100	a=893827;b=-419296;opcode=000;
			#100	a=547627;b=193168;opcode=100;
			#100	a=57904;b=-539019;opcode=111;
			#100	a=-197922;b=-290877;opcode=010;
			#100	a=-281373;b=-576893;opcode=110;
			#100	a=-198299;b=529217;opcode=010;
			#100	a=-865885;b=854955;opcode=000;
			#100	a=683892;b=685561;opcode=001;
			#100	a=90427;b=383451;opcode=000;
			#100	a=-970443;b=105955;opcode=111;
			#100	a=250382;b=890409;opcode=000;
			#100	a=494244;b=-553912;opcode=100;
			#100	a=844009;b=-15147;opcode=110;
			#100	a=134343;b=910540;opcode=111;
			#100	a=655089;b=145791;opcode=010;
			#100	a=335469;b=-519475;opcode=001;
			#100	a=-388294;b=-151552;opcode=111;
			#100	a=-754682;b=-813605;opcode=010;
			#100	a=431647;b=795051;opcode=110;
			#100	a=141497;b=773488;opcode=100;
			#100	a=-588127;b=-641422;opcode=001;
			#100	a=-918968;b=10109;opcode=001;
			#100	a=710850;b=584937;opcode=000;
			#100	a=-419276;b=-931897;opcode=010;
			#100	a=499616;b=230242;opcode=001;
			#100	a=-598168;b=-515282;opcode=010;
			#100	a=509327;b=-750238;opcode=010;
			#100	a=-345293;b=-695833;opcode=100;
			#100	a=99982;b=809622;opcode=000;
			#100	a=-994158;b=-503542;opcode=100;
			#100	a=552661;b=671341;opcode=000;
			#100	a=-791722;b=690684;opcode=000;
			#100	a=-11136;b=785467;opcode=001;
			#100	a=547280;b=37907;opcode=001;
			#100	a=-180054;b=-941005;opcode=111;
			#100	a=-957327;b=347129;opcode=001;
			#100	a=401421;b=530612;opcode=110;
			#100	a=-186477;b=-957005;opcode=010;
			#100	a=60260;b=-810816;opcode=100;
			#100	a=578062;b=246251;opcode=110;
			#100	a=-825161;b=-859572;opcode=111;
			#100	a=24488;b=-50280;opcode=110;
			#100	a=636129;b=287941;opcode=000;
			#100	a=-170033;b=739547;opcode=010;
			#100	a=5505;b=-771421;opcode=110;
			#100	a=-812407;b=713635;opcode=110;
			#100	a=110088;b=874031;opcode=100;
			#100	a=877531;b=325391;opcode=110;
			#100	a=917726;b=696056;opcode=111;
			#100	a=312458;b=-618468;opcode=001;
			#100	a=111071;b=850460;opcode=111;
			#100	a=-503091;b=-761734;opcode=010;
			#100	a=365010;b=169873;opcode=110;
			#100	a=1522;b=541130;opcode=110;
			#100	a=258431;b=-478334;opcode=001;
			#100	a=369223;b=-375073;opcode=100;
			#100	a=-405045;b=641079;opcode=110;
			#100	a=-818163;b=-816134;opcode=001;
			#100	a=590411;b=-96923;opcode=100;
			#100	a=-648892;b=-630021;opcode=000;
			#100	a=56076;b=233841;opcode=001;
			#100	a=857625;b=371080;opcode=110;
			#100	a=805436;b=762983;opcode=100;
			#100	a=951844;b=156816;opcode=111;
			#100	a=-342407;b=865042;opcode=111;
			#100	a=313175;b=835737;opcode=111;
			#100	a=-786144;b=405162;opcode=001;
			#100	a=163564;b=257298;opcode=001;
			#100	a=615127;b=611122;opcode=110;
			#100	a=-952338;b=977028;opcode=111;
			#100	a=-981;b=495837;opcode=110;
			#100	a=454238;b=-786072;opcode=100;
			#100	a=628822;b=-313677;opcode=111;
			#100	a=269302;b=556827;opcode=010;
			#100	a=-150999;b=-900192;opcode=100;
			#100	a=-578278;b=-736821;opcode=010;
			#100	a=350717;b=666056;opcode=110;
			#100	a=45401;b=878041;opcode=001;
			#100	a=-975793;b=-572137;opcode=111;
			#100	a=684488;b=-24526;opcode=001;
			#100	a=243595;b=837900;opcode=000;
			#100	a=183887;b=-382133;opcode=001;
			#100	a=-33431;b=-743749;opcode=001;
			#100	a=-869646;b=-998099;opcode=110;
			#100	a=-98021;b=-498768;opcode=001;
			#100	a=235417;b=-283463;opcode=100;
			#100	a=555975;b=554562;opcode=001;
			#100	a=937410;b=19230;opcode=010;
			#100	a=-441057;b=926069;opcode=010;
			#100	a=-607382;b=-463850;opcode=000;
			#100	a=-289077;b=240140;opcode=110;
			#100	a=316105;b=302448;opcode=010;
			#100	a=-98597;b=842292;opcode=010;
			#100	a=550300;b=937315;opcode=001;
			#100	a=407626;b=-838191;opcode=100;
			#100	a=-219091;b=-460096;opcode=111;
			#100	a=-96025;b=127844;opcode=111;
			#100	a=47525;b=144965;opcode=001;
			#100	a=535889;b=777515;opcode=110;
			#100	a=-566476;b=-7541;opcode=110;
			#100	a=-274967;b=-798915;opcode=110;
			#100	a=-933374;b=-22618;opcode=010;
			#100	a=-590967;b=-230735;opcode=111;
			#100	a=242130;b=-921224;opcode=100;
			#100	a=537398;b=-28467;opcode=010;
			#100	a=358399;b=-620068;opcode=100;
			#100	a=-731407;b=542626;opcode=100;
			#100	a=652312;b=745129;opcode=000;
			#100	a=-327647;b=889511;opcode=100;
			#100	a=-956705;b=-997757;opcode=010;
			#100	a=930671;b=-235378;opcode=110;
			#100	a=-260639;b=472897;opcode=111;
			#100	a=-625480;b=808424;opcode=000;
			#100	a=-460026;b=872892;opcode=000;
			#100	a=404849;b=897901;opcode=000;
			#100	a=865340;b=866085;opcode=110;
			#100	a=569548;b=-154556;opcode=100;
			#100	a=135880;b=-114553;opcode=010;
			#100	a=-777907;b=-59692;opcode=000;
			#100	a=434956;b=713185;opcode=010;
			#100	a=-205638;b=-6867;opcode=010;
			#100	a=-806009;b=-107689;opcode=111;
			#100	a=564091;b=590848;opcode=010;
			#100	a=340847;b=913499;opcode=010;
			#100	a=-901750;b=-849706;opcode=111;
			#100	a=278504;b=-828441;opcode=001;
			#100	a=-675751;b=734797;opcode=100;
			#100	a=-239095;b=54353;opcode=111;
			#100	a=-142000;b=466369;opcode=110;
			#100	a=699461;b=566034;opcode=010;
			#100	a=781812;b=-144873;opcode=001;
			#100	a=-732358;b=309820;opcode=010;
			#100	a=776111;b=-207998;opcode=000;
			#100	a=-461940;b=893082;opcode=100;
			#100	a=-579114;b=590933;opcode=010;
			#100	a=568295;b=-672911;opcode=001;
			#100	a=-312808;b=516162;opcode=000;
			#100	a=-164858;b=595106;opcode=001;
			#100	a=-727800;b=875700;opcode=110;
			#100	a=593213;b=571617;opcode=110;
			#100	a=-949266;b=-488623;opcode=001;
			#100	a=974526;b=672677;opcode=110;
			#100	a=254661;b=-841333;opcode=000;
			#100	a=-140226;b=279833;opcode=110;
			#100	a=796785;b=-799854;opcode=110;
			#100	a=-607747;b=-361075;opcode=010;
			#100	a=186202;b=105915;opcode=001;
			#100	a=82004;b=105112;opcode=001;
			#100	a=-474307;b=-481568;opcode=110;
			#100	a=-230262;b=745346;opcode=001;
			#100	a=-840951;b=-932187;opcode=111;
			#100	a=-813749;b=-244653;opcode=010;
			#100	a=-629949;b=-130001;opcode=100;
			#100	a=802816;b=-734452;opcode=001;
			#100	a=-759168;b=788372;opcode=001;
			#100	a=513008;b=-177525;opcode=100;
			#100	a=-81920;b=20382;opcode=010;
			#100	a=144157;b=-760453;opcode=001;
			#100	a=-123062;b=-779015;opcode=001;
			#100	a=-705603;b=-331785;opcode=001;
			#100	a=521000;b=-550468;opcode=100;
			#100	a=943176;b=346040;opcode=100;
			#100	a=163494;b=517981;opcode=110;
			#100	a=78782;b=86411;opcode=010;
			#100	a=906211;b=-981678;opcode=001;
			#100	a=283887;b=635365;opcode=100;
			#100	a=-609821;b=-987014;opcode=111;
			#100	a=498180;b=-408565;opcode=100;
			#100	a=-669536;b=-961008;opcode=110;
			#100	a=296926;b=-677857;opcode=000;
			#100	a=-992501;b=-126237;opcode=010;
			#100	a=-115485;b=-95235;opcode=001;
			#100	a=795643;b=237373;opcode=110;
			#100	a=-87168;b=210344;opcode=010;
			#100	a=-605281;b=-683003;opcode=000;
			#100	a=-714285;b=-333444;opcode=001;
			#100	a=358578;b=995764;opcode=000;
			#100	a=-658179;b=258290;opcode=001;
			#100	a=-230218;b=-766173;opcode=111;
			#100	a=-182557;b=30601;opcode=111;
			#100	a=531870;b=935749;opcode=110;
			#100	a=464716;b=-870925;opcode=010;
			#100	a=887538;b=140620;opcode=100;
			#100	a=642404;b=145703;opcode=111;
			#100	a=685314;b=109890;opcode=100;
			#100	a=-189169;b=87143;opcode=010;
			#100	a=-450430;b=384492;opcode=100;
			#100	a=-23106;b=564786;opcode=001;
			#100	a=-922308;b=-790126;opcode=000;
			#100	a=-264920;b=-258534;opcode=110;
			#100	a=-533083;b=-270529;opcode=010;
			#100	a=860255;b=-435894;opcode=111;
			#100	a=-108814;b=-499146;opcode=110;
			#100	a=301236;b=-910675;opcode=001;
			#100	a=733834;b=-349871;opcode=010;
			#100	a=919327;b=811155;opcode=110;
			#100	a=324719;b=6991;opcode=010;
			#100	a=836241;b=693061;opcode=000;
			#100	a=113245;b=-964364;opcode=010;
			#100	a=-544815;b=-214348;opcode=010;
			#100	a=-622863;b=540020;opcode=001;
			#100	a=-297678;b=114110;opcode=110;
			#100	a=706152;b=271007;opcode=111;
			#100	a=443612;b=-382926;opcode=010;
			#100	a=776619;b=-6085;opcode=111;
			#100	a=457615;b=920070;opcode=001;
			#100	a=-182496;b=541358;opcode=111;
			#100	a=340834;b=-827078;opcode=000;
			#100	a=769570;b=125129;opcode=010;
			#100	a=735477;b=-56300;opcode=001;
			#100	a=-272543;b=-623749;opcode=010;
			#100	a=-749711;b=582674;opcode=100;
			#100	a=-624691;b=380205;opcode=111;
			#100	a=833341;b=-8238;opcode=110;
			#100	a=216558;b=-538497;opcode=100;
			#100	a=-478702;b=-62791;opcode=010;
			#100	a=-235230;b=600854;opcode=110;
			#100	a=334280;b=-105420;opcode=100;
			#100	a=-289985;b=210093;opcode=100;
			#100	a=-567124;b=-849546;opcode=000;
			#100	a=225872;b=221319;opcode=100;
			#100	a=-102948;b=601359;opcode=010;
			#100	a=176641;b=467493;opcode=000;
			#100	a=421432;b=-122476;opcode=111;
			#100	a=-375007;b=36851;opcode=111;
			#100	a=-433478;b=-734683;opcode=100;
			#100	a=55055;b=-127476;opcode=100;
			#100	a=-84416;b=848349;opcode=000;
			#100	a=-499509;b=603554;opcode=111;
			#100	a=736451;b=-331855;opcode=001;
			#100	a=423008;b=-42221;opcode=010;
			#100	a=-537876;b=-613202;opcode=001;
			#100	a=902865;b=-864200;opcode=001;
			#100	a=-308696;b=-491217;opcode=001;
			#100	a=-581323;b=597703;opcode=010;
			#100	a=349037;b=-39119;opcode=100;
			#100	a=828889;b=69443;opcode=001;
			#100	a=-724554;b=238129;opcode=000;
			#100	a=127322;b=-813953;opcode=110;
			#100	a=-334078;b=723648;opcode=100;
			#100	a=-543054;b=824879;opcode=100;
			#100	a=-381554;b=154474;opcode=110;
			#100	a=421223;b=176912;opcode=111;
			#100	a=69699;b=-44924;opcode=111;
			#100	a=39727;b=-860155;opcode=000;
			#100	a=-340602;b=-233212;opcode=001;
			#100	a=361191;b=-965414;opcode=111;
			#100	a=786602;b=-417285;opcode=010;
			#100	a=-309271;b=-982052;opcode=110;
			#100	a=-305155;b=124562;opcode=010;
			#100	a=662934;b=-331881;opcode=110;
			#100	a=332406;b=-55319;opcode=001;
			#100	a=135801;b=-141630;opcode=010;
			#100	a=660526;b=-133772;opcode=100;
			#100	a=-534665;b=-102994;opcode=010;
			#100	a=33975;b=98218;opcode=100;
			#100	a=971370;b=-263491;opcode=110;
			#100	a=-365721;b=921231;opcode=010;
			#100	a=140105;b=-820994;opcode=001;
			#100	a=217425;b=-253160;opcode=111;
			#100	a=194150;b=519977;opcode=111;
			#100	a=684087;b=155275;opcode=110;
			#100	a=-710295;b=511961;opcode=000;
			#100	a=27992;b=-824404;opcode=010;
			#100	a=-828925;b=380092;opcode=000;
			#100	a=-484431;b=252285;opcode=111;
			#100	a=-657851;b=-516928;opcode=111;
			#100	a=864308;b=640311;opcode=110;
			#100	a=684350;b=-305206;opcode=001;
			#100	a=164390;b=370096;opcode=000;
			#100	a=96581;b=-474027;opcode=110;
			#100	a=-742190;b=-718809;opcode=010;
			#100	a=-668769;b=-924637;opcode=001;
			#100	a=712032;b=943021;opcode=111;
			#100	a=132385;b=-637763;opcode=010;
			#100	a=-80800;b=888777;opcode=111;
			#100	a=-470832;b=677768;opcode=010;
			#100	a=166883;b=-798735;opcode=010;
			#100	a=-776454;b=371415;opcode=010;
			#100	a=583980;b=-334585;opcode=110;
			#100	a=-148473;b=477839;opcode=110;
			#100	a=-344697;b=654900;opcode=000;
			#100	a=-370715;b=-172137;opcode=000;
			#100	a=-638391;b=935693;opcode=010;
			#100	a=209744;b=-649910;opcode=110;
			#100	a=-192113;b=-273717;opcode=110;
			#100	a=958;b=-504741;opcode=000;
			#100	a=-932504;b=972002;opcode=111;
			#100	a=-426347;b=-212083;opcode=110;
			#100	a=-14153;b=-751947;opcode=001;
			#100	a=-430216;b=561864;opcode=110;
			#100	a=928302;b=-656531;opcode=010;
			#100	a=738487;b=942828;opcode=001;
			#100	a=885786;b=-835481;opcode=110;
			#100	a=-628660;b=242632;opcode=110;
			#100	a=339560;b=-963441;opcode=100;
			#100	a=508450;b=683497;opcode=111;
			#100	a=991080;b=698118;opcode=100;
			#100	a=-396956;b=-596464;opcode=010;
			#100	a=468311;b=880095;opcode=001;
			#100	a=736140;b=102089;opcode=000;
			#100	a=763037;b=491849;opcode=100;
			#100	a=-920792;b=755404;opcode=100;
			#100	a=-447246;b=-521850;opcode=100;
			#100	a=-630490;b=425839;opcode=001;
			#100	a=-9261;b=-665108;opcode=111;
			#100	a=599055;b=499286;opcode=010;
			#100	a=310523;b=-60589;opcode=000;
			#100	a=794032;b=146253;opcode=110;
			#100	a=737946;b=995600;opcode=100;
			#100	a=892770;b=-608442;opcode=100;
			#100	a=857217;b=-598645;opcode=110;
			#100	a=876130;b=842142;opcode=001;
			#100	a=616466;b=551245;opcode=000;
			#100	a=547843;b=668250;opcode=001;
			#100	a=150248;b=-619462;opcode=111;
			#100	a=-992582;b=937335;opcode=110;
			#100	a=256268;b=399862;opcode=001;
			#100	a=-785799;b=-566098;opcode=110;
			#100	a=167884;b=-309159;opcode=000;
			#100	a=980738;b=989031;opcode=111;
			#100	a=250532;b=-25309;opcode=000;
			#100	a=43812;b=486193;opcode=110;
			#100	a=36762;b=453410;opcode=100;
			#100	a=-677282;b=366452;opcode=111;
			#100	a=-423675;b=313645;opcode=001;
			#100	a=807184;b=798793;opcode=111;
			#100	a=-64479;b=-14520;opcode=000;
			#100	a=-105701;b=-222018;opcode=001;
			#100	a=-131995;b=-781802;opcode=110;
			#100	a=-834399;b=212087;opcode=010;
			#100	a=335418;b=-18044;opcode=010;
			#100	a=117507;b=-669063;opcode=100;
			#100	a=-202892;b=531839;opcode=110;
			#100	a=-397580;b=950459;opcode=110;
			#100	a=-57053;b=210173;opcode=000;
			#100	a=-877762;b=929740;opcode=100;
			#100	a=174237;b=832683;opcode=111;
			#100	a=82210;b=-126546;opcode=001;
			#100	a=-636201;b=-606108;opcode=001;
			#100	a=139427;b=879626;opcode=110;
			#100	a=825280;b=91118;opcode=001;
			#100	a=246948;b=464055;opcode=010;
			#100	a=-462544;b=112367;opcode=010;
			#100	a=-886294;b=223570;opcode=111;
			#100	a=-335725;b=650516;opcode=100;
			#100	a=909210;b=10293;opcode=001;
			#100	a=-701359;b=369788;opcode=000;
			#100	a=-863538;b=397208;opcode=100;
			#100	a=867140;b=179669;opcode=010;
			#100	a=918205;b=-314490;opcode=000;
			#100	a=340098;b=591589;opcode=100;
			#100	a=365928;b=8330;opcode=111;
			#100	a=341984;b=-54052;opcode=010;
			#100	a=-755675;b=-388377;opcode=010;
			#100	a=195980;b=-357285;opcode=100;
			#100	a=934112;b=-435486;opcode=000;
			#100	a=-547568;b=-663155;opcode=010;
			#100	a=-718644;b=-29435;opcode=001;
			#100	a=-537647;b=-589340;opcode=111;
			#100	a=-150648;b=-638226;opcode=010;
			#100	a=405189;b=731203;opcode=111;
			#100	a=178064;b=-608768;opcode=110;
			#100	a=872832;b=277194;opcode=100;
			#100	a=-153295;b=990712;opcode=111;
			#100	a=196518;b=73966;opcode=100;
			#100	a=496709;b=340136;opcode=100;
			#100	a=294410;b=-238091;opcode=110;
			#100	a=-755946;b=-674921;opcode=110;
			#100	a=-400957;b=-448490;opcode=010;
			#100	a=-519486;b=-528777;opcode=001;
			#100	a=327741;b=-414298;opcode=001;
			#100	a=-470088;b=860769;opcode=010;
			#100	a=-349566;b=-779668;opcode=010;
			#100	a=218639;b=-132490;opcode=111;
			#100	a=89733;b=543355;opcode=010;
			#100	a=580840;b=-396957;opcode=001;
			#100	a=-291846;b=-713593;opcode=111;
			#100	a=-921953;b=-776452;opcode=111;
			#100	a=687246;b=557400;opcode=110;
			#100	a=31666;b=-168076;opcode=010;
			#100	a=-882212;b=758266;opcode=000;
			#100	a=795394;b=-861567;opcode=000;
			#100	a=702711;b=720882;opcode=010;
			#100	a=-14013;b=-570579;opcode=110;
			#100	a=-887939;b=-237113;opcode=110;
			#100	a=-574402;b=482267;opcode=100;
			#100	a=386246;b=151124;opcode=000;
			#100	a=193195;b=987788;opcode=010;
			#100	a=-838450;b=726800;opcode=000;
			#100	a=473574;b=-37219;opcode=001;
			#100	a=-275088;b=119228;opcode=110;
			#100	a=-952209;b=118466;opcode=000;
			#100	a=-239962;b=526279;opcode=001;
			#100	a=809336;b=333819;opcode=110;
			#100	a=249244;b=430771;opcode=100;
			#100	a=-331805;b=962005;opcode=001;
			#100	a=34029;b=-550438;opcode=110;
			#100	a=561576;b=-381768;opcode=000;
			#100	a=-960151;b=-327474;opcode=111;
			#100	a=-367223;b=-477470;opcode=111;
			#100	a=-726786;b=-706147;opcode=001;
			#100	a=-374225;b=-301370;opcode=000;
			#100	a=-709822;b=979467;opcode=001;
			#100	a=-168870;b=-251945;opcode=111;
			#100	a=-795588;b=955094;opcode=000;
			#100	a=850970;b=-592883;opcode=001;
			#100	a=-447644;b=55177;opcode=010;
			#100	a=-733226;b=-471690;opcode=010;
			#100	a=17198;b=426785;opcode=010;
			#100	a=732937;b=390699;opcode=000;
			#100	a=377636;b=772992;opcode=110;
			#100	a=17342;b=-464588;opcode=111;
			#100	a=417648;b=887125;opcode=000;
			#100	a=-257468;b=545102;opcode=000;
			#100	a=-894719;b=-264047;opcode=000;
			#100	a=346864;b=-650399;opcode=001;
			#100	a=-160441;b=-661384;opcode=001;
			#100	a=125463;b=-981673;opcode=001;
			#100	a=792566;b=299716;opcode=110;
			#100	a=-137209;b=975014;opcode=100;
			#100	a=962148;b=925322;opcode=100;
			#100	a=78053;b=670585;opcode=100;
			#100	a=-354588;b=-504810;opcode=000;
			#100	a=-488588;b=-467266;opcode=010;
			#100	a=-222392;b=347195;opcode=000;
			#100	a=-52483;b=317246;opcode=110;
			#100	a=564368;b=770324;opcode=001;
			#100	a=-977819;b=-168437;opcode=010;
			#100	a=809674;b=676796;opcode=100;
			#100	a=699177;b=-602035;opcode=001;
			#100	a=262449;b=-760349;opcode=010;
			#100	a=323570;b=-973321;opcode=000;
			#100	a=-77188;b=30563;opcode=001;
			#100	a=915654;b=-870599;opcode=010;
			#100	a=474168;b=-360062;opcode=010;
			#100	a=129881;b=-260791;opcode=100;
			#100	a=387165;b=-315086;opcode=110;
			#100	a=623730;b=359011;opcode=110;
			#100	a=57705;b=-800016;opcode=001;
			#100	a=-883663;b=830473;opcode=111;
			#100	a=-357297;b=462973;opcode=000;
			#100	a=176405;b=739313;opcode=110;
			#100	a=-719237;b=61430;opcode=000;
			#100	a=-197159;b=-490697;opcode=000;
			#100	a=-541812;b=719528;opcode=100;
			#100	a=802977;b=328335;opcode=110;
			#100	a=709863;b=822122;opcode=110;
			#100	a=320254;b=51117;opcode=100;
			#100	a=736316;b=818742;opcode=110;
			#100	a=-611600;b=139649;opcode=001;
			#100	a=-659024;b=-228041;opcode=111;
			#100	a=-539181;b=-561745;opcode=111;
			#100	a=827175;b=983961;opcode=000;
			#100	a=-808787;b=276686;opcode=001;
			#100	a=446525;b=602315;opcode=100;
			#100	a=-395977;b=-473178;opcode=111;
			#100	a=-309065;b=-517901;opcode=111;
			#100	a=529027;b=-965463;opcode=001;
			#100	a=23872;b=424457;opcode=000;
			#100	a=-1235;b=226585;opcode=001;
			#100	a=615375;b=-829017;opcode=110;
			#100	a=-748524;b=570675;opcode=001;
			#100	a=-380640;b=-742615;opcode=100;
			#100	a=314685;b=340448;opcode=001;
			#100	a=-147819;b=-48177;opcode=100;
			#100	a=999991;b=988728;opcode=110;
			#100	a=394483;b=-368694;opcode=111;
			#100	a=-41790;b=-982221;opcode=010;
			#100	a=-951225;b=-217313;opcode=000;
			#100	a=-944143;b=-349350;opcode=000;
			#100	a=-927183;b=148920;opcode=001;
			#100	a=-690276;b=650890;opcode=001;
			#100	a=698107;b=993350;opcode=000;
			#100	a=284384;b=-598967;opcode=001;
			#100	a=-372088;b=-141552;opcode=110;
			#100	a=712684;b=363890;opcode=100;
			#100	a=-332806;b=-852235;opcode=000;
			#100	a=-225748;b=-522008;opcode=000;
			#100	a=-932378;b=-702678;opcode=110;
			#100	a=-772308;b=443239;opcode=001;
			#100	a=-901715;b=169377;opcode=000;
			#100	a=-294965;b=812176;opcode=010;
			#100	a=-358340;b=-68710;opcode=001;
			#100	a=800356;b=-223269;opcode=000;
			#100	a=183613;b=-447770;opcode=000;
			#100	a=-363362;b=-949370;opcode=111;
			#100	a=-754471;b=-824001;opcode=000;
			#100	a=740459;b=115313;opcode=110;
			#100	a=680714;b=792611;opcode=001;
			#100	a=608495;b=185601;opcode=000;
			#100	a=-254707;b=995652;opcode=100;
			#100	a=-656240;b=-182244;opcode=001;
			#100	a=581713;b=915874;opcode=111;
			#100	a=-142651;b=-655820;opcode=110;
			#100	a=265693;b=-775047;opcode=110;
			#100	a=409561;b=-722845;opcode=100;
			#100	a=-385460;b=589049;opcode=001;
			#100	a=-836944;b=-213916;opcode=111;
			#100	a=663191;b=-323143;opcode=000;
			#100	a=772526;b=-949687;opcode=010;
			#100	a=419054;b=848051;opcode=110;
			#100	a=556881;b=-474764;opcode=010;
			#100	a=8432;b=437173;opcode=001;
			#100	a=52189;b=-127147;opcode=000;
			#100	a=-632842;b=803392;opcode=000;
			#100	a=-457806;b=-259713;opcode=110;
			#100	a=-927856;b=303621;opcode=001;
			#100	a=481987;b=917147;opcode=001;
			#100	a=1682;b=-227134;opcode=110;
			#100	a=-584719;b=-730533;opcode=001;
			#100	a=-390207;b=879360;opcode=001;
			#100	a=315625;b=-313677;opcode=001;
			#100	a=-637332;b=508978;opcode=110;
			#100	a=746282;b=-505489;opcode=001;
			#100	a=-813920;b=-39932;opcode=110;
			#100	a=-212166;b=116222;opcode=010;
			#100	a=-624514;b=944377;opcode=100;
			#100	a=183598;b=202516;opcode=111;
			#100	a=266694;b=591385;opcode=010;
			#100	a=-313300;b=900604;opcode=001;
			#100	a=-876439;b=-300914;opcode=110;
			#100	a=437100;b=392050;opcode=010;
			#100	a=-204491;b=-631698;opcode=110;
			#100	a=-611557;b=-20477;opcode=110;
			#100	a=-459844;b=-15262;opcode=000;
			#100	a=-419580;b=987213;opcode=001;
			#100	a=-275482;b=197678;opcode=111;
			#100	a=-464338;b=-829921;opcode=100;
			#100	a=941628;b=-628313;opcode=010;
			#100	a=-831323;b=211163;opcode=110;
			#100	a=610777;b=-56846;opcode=001;
			#100	a=-22033;b=452166;opcode=100;
			#100	a=-81273;b=-273271;opcode=100;
			#100	a=-266472;b=403005;opcode=010;
			#100	a=-44150;b=-784136;opcode=110;
			#100	a=-742916;b=113704;opcode=000;
			#100	a=840508;b=181911;opcode=010;
			#100	a=-918590;b=212992;opcode=010;
			#100	a=-724239;b=-800463;opcode=110;
			#100	a=-794665;b=-215791;opcode=100;
			#100	a=-768735;b=705058;opcode=001;
			#100	a=-348313;b=-247527;opcode=100;
			#100	a=-886161;b=-425184;opcode=010;
			#100	a=-915698;b=-958850;opcode=010;
			#100	a=-965865;b=-878549;opcode=100;
			#100	a=-373084;b=927725;opcode=111;
			#100	a=468204;b=595277;opcode=111;
			#100	a=-867138;b=357576;opcode=111;
			#100	a=-528197;b=913386;opcode=100;
			#100	a=879955;b=185172;opcode=111;
			#100	a=-151857;b=-226573;opcode=100;
			#100	a=476158;b=458242;opcode=001;
			#100	a=111232;b=818722;opcode=111;
			#100	a=185133;b=-89399;opcode=000;
			#100	a=-319422;b=-871421;opcode=111;
			#100	a=-244360;b=-448393;opcode=111;
			#100	a=-334936;b=-9485;opcode=110;
			#100	a=-959430;b=-210211;opcode=010;
			#100	a=-104796;b=-446934;opcode=001;
			#100	a=788131;b=113780;opcode=001;
			#100	a=-945782;b=777367;opcode=100;
			#100	a=-274339;b=648340;opcode=000;
			#100	a=-503291;b=-371090;opcode=110;
			#100	a=-754542;b=372879;opcode=110;
			#100	a=-289421;b=-285683;opcode=001;
			#100	a=576631;b=516308;opcode=110;
			#100	a=307232;b=298906;opcode=110;
			#100	a=426831;b=239292;opcode=010;
			#100	a=283012;b=769539;opcode=000;
			#100	a=147508;b=668596;opcode=001;
			#100	a=394607;b=-65659;opcode=000;
			#100	a=644020;b=925578;opcode=110;
			#100	a=827629;b=-940561;opcode=111;
			#100	a=374547;b=-999765;opcode=111;
			#100	a=69508;b=-82089;opcode=010;
			#100	a=-512721;b=-446117;opcode=110;
			#100	a=143411;b=506891;opcode=110;
			#100	a=175239;b=-210525;opcode=001;
			#100	a=727730;b=-65187;opcode=000;
			#100	a=-950201;b=-379860;opcode=111;
			#100	a=358768;b=-831731;opcode=010;
			#100	a=-309804;b=-612600;opcode=010;
			#100	a=812825;b=-115212;opcode=010;
			#100	a=438178;b=-173316;opcode=000;
			#100	a=552695;b=-631090;opcode=111;
			#100	a=-535716;b=-964319;opcode=111;
			#100	a=-962640;b=-642809;opcode=001;
			#100	a=690326;b=289014;opcode=110;
			#100	a=-312531;b=-358680;opcode=111;
			#100	a=-575;b=-451280;opcode=100;
			#100	a=930193;b=-698191;opcode=001;
			#100	a=348204;b=-508614;opcode=010;
			#100	a=-5024;b=91765;opcode=110;
			#100	a=335453;b=-177550;opcode=110;
			#100	a=673083;b=740761;opcode=000;
			#100	a=-32214;b=984539;opcode=000;
			#100	a=802800;b=453244;opcode=000;
			#100	a=-54396;b=166306;opcode=111;
			#100	a=-310120;b=462320;opcode=100;
			#100	a=-349033;b=836756;opcode=000;
			#100	a=-283791;b=444781;opcode=001;
			#100	a=-840246;b=333718;opcode=010;
			#100	a=34580;b=-995194;opcode=111;
			#100	a=-369145;b=381165;opcode=110;
			#100	a=360574;b=-759961;opcode=111;
			#100	a=-12367;b=-262460;opcode=000;
			#100	a=90367;b=802378;opcode=111;
			#100	a=795608;b=-256436;opcode=100;
			#100	a=-503958;b=436039;opcode=111;
			#100	a=-556283;b=10834;opcode=000;
			#100	a=-802995;b=325642;opcode=100;
			#100	a=-701366;b=736342;opcode=110;
			#100	a=910985;b=304142;opcode=100;
			#100	a=-530369;b=-790994;opcode=100;
			#100	a=-397297;b=-801336;opcode=001;
			#100	a=689253;b=-795538;opcode=000;
			#100	a=926365;b=978342;opcode=010;
			#100	a=261205;b=5655;opcode=110;
			#100	a=122281;b=334934;opcode=000;
			#100	a=988002;b=-103498;opcode=000;
			#100	a=-455821;b=-353615;opcode=100;
			#100	a=-798479;b=8297;opcode=110;
			#100	a=416370;b=591726;opcode=110;
			#100	a=-989767;b=-227767;opcode=100;
			#100	a=-298703;b=799085;opcode=010;
			#100	a=-718020;b=-887382;opcode=100;
			#100	a=197777;b=-801514;opcode=110;
			#100	a=192931;b=-411740;opcode=000;
			#100	a=519930;b=238446;opcode=111;
			#100	a=124538;b=-550239;opcode=001;
			#100	a=-692207;b=408488;opcode=111;
			#100	a=39803;b=-159158;opcode=000;
			#100	a=392957;b=394310;opcode=000;
			#100	a=686663;b=265039;opcode=000;
			#100	a=-137686;b=-773222;opcode=100;
			#100	a=250578;b=-634570;opcode=010;
			#100	a=-97354;b=850564;opcode=111;
			#100	a=841429;b=-282841;opcode=010;
			#100	a=564198;b=-170600;opcode=110;
			#100	a=962624;b=-308909;opcode=010;
			#100	a=778977;b=743670;opcode=001;
			#100	a=-989508;b=-350014;opcode=111;
			#100	a=575076;b=-283394;opcode=100;
			#100	a=-960159;b=396324;opcode=111;
			#100	a=-959771;b=-488505;opcode=000;
			#100	a=886034;b=839671;opcode=001;
			#100	a=-80207;b=-960580;opcode=010;
			#100	a=671178;b=108124;opcode=010;
			#100	a=482151;b=195656;opcode=100;
			#100	a=-59973;b=-249710;opcode=000;
			#100	a=-741315;b=786976;opcode=001;
			#100	a=340796;b=-965824;opcode=110;
			#100	a=857404;b=592364;opcode=100;
			#100	a=-223016;b=394026;opcode=001;
			#100	a=-301692;b=51214;opcode=110;
			#100	a=416599;b=-836559;opcode=111;
			#100	a=-634610;b=-421350;opcode=001;
			#100	a=-187047;b=-185693;opcode=111;
			#100	a=-56495;b=-953614;opcode=100;
			#100	a=-194643;b=-290879;opcode=110;
			#100	a=-532162;b=454779;opcode=000;
			#100	a=87709;b=-618402;opcode=001;
			#100	a=313078;b=356577;opcode=110;
			#100	a=-974649;b=-263662;opcode=111;
			#100	a=115902;b=12376;opcode=111;
			#100	a=-216095;b=-903546;opcode=111;
			#100	a=-184468;b=-147944;opcode=001;
			#100	a=250668;b=515357;opcode=100;
			#100	a=-177119;b=-975579;opcode=010;
			#100	a=243411;b=55744;opcode=111;
			#100	a=-831148;b=164208;opcode=001;
			#100	a=511218;b=-569400;opcode=010;
			#100	a=853450;b=275441;opcode=001;
			#100	a=-449682;b=197375;opcode=001;
			#100	a=-492491;b=538200;opcode=110;
			#100	a=209812;b=486748;opcode=001;
			#100	a=-287326;b=280257;opcode=110;
			#100	a=-851212;b=-148851;opcode=110;
			#100	a=294587;b=753558;opcode=111;
			#100	a=-486818;b=-212591;opcode=110;
			#100	a=-861353;b=-164217;opcode=111;
			#100	a=-238070;b=-409635;opcode=001;
			#100	a=-520804;b=66912;opcode=000;
			#100	a=-378131;b=550834;opcode=111;
			#100	a=-561176;b=-4254;opcode=100;
			#100	a=804503;b=-546753;opcode=001;
			#100	a=890901;b=542318;opcode=001;
			#100	a=895558;b=-441596;opcode=100;
			#100	a=-397925;b=597647;opcode=110;
			#100	a=443355;b=146756;opcode=010;
			#100	a=179794;b=307863;opcode=010;
			#100	a=222453;b=-103014;opcode=100;
			#100	a=-537397;b=-448345;opcode=100;
			#100	a=-140307;b=30074;opcode=111;
			#100	a=-413192;b=385933;opcode=010;
			#100	a=818237;b=377212;opcode=100;
			#100	a=729026;b=-294786;opcode=000;
			#100	a=715480;b=980667;opcode=001;
			#100	a=120499;b=-90844;opcode=000;
			#100	a=-988813;b=541518;opcode=001;
			#100	a=978995;b=-246269;opcode=001;
			#100	a=-39161;b=127897;opcode=110;
			#100	a=-995270;b=637089;opcode=111;
			#100	a=134903;b=322582;opcode=001;
			#100	a=396304;b=218474;opcode=010;
			#100	a=-747502;b=-560872;opcode=110;
			#100	a=586853;b=-890983;opcode=100;
			#100	a=898345;b=-706179;opcode=000;
			#100	a=419173;b=-72750;opcode=100;
			#100	a=235068;b=-570376;opcode=100;
			#100	a=-468565;b=-564067;opcode=000;
			#100	a=-414136;b=-472675;opcode=110;
			#100	a=-161710;b=840206;opcode=111;
			#100	a=689904;b=-42336;opcode=001;
			#100	a=153723;b=-979781;opcode=110;
			#100	a=-285021;b=265697;opcode=001;
			#100	a=336077;b=463764;opcode=100;
			#100	a=333803;b=519338;opcode=111;
			#100	a=-623165;b=-446841;opcode=001;
			#100	a=242516;b=184236;opcode=001;
			#100	a=158196;b=-730836;opcode=001;
			#100	a=-362359;b=826158;opcode=000;
			#100	a=-168854;b=199634;opcode=110;
			#100	a=-508051;b=817536;opcode=001;
			#100	a=578071;b=-276637;opcode=111;
			#100	a=-210853;b=888323;opcode=000;
			#100	a=-692714;b=-162090;opcode=100;
			#100	a=-604422;b=-140769;opcode=110;
			#100	a=697003;b=-404940;opcode=010;
			#100	a=-319621;b=-742130;opcode=000;
			#100	a=906915;b=451953;opcode=010;
			#100	a=-40919;b=438743;opcode=001;
			#100	a=659114;b=-33366;opcode=111;
			#100	a=-539811;b=529134;opcode=110;
			#100	a=812615;b=204526;opcode=111;
			#100	a=-475977;b=-250268;opcode=010;
			#100	a=-273129;b=166809;opcode=010;
			#100	a=-212206;b=-203190;opcode=010;
			#100	a=-429872;b=223594;opcode=111;
			#100	a=672013;b=-144279;opcode=100;
			#100	a=-658059;b=640613;opcode=001;
			#100	a=644502;b=419522;opcode=001;
			#100	a=738139;b=-847118;opcode=000;
			#100	a=-530786;b=-665662;opcode=111;
			#100	a=-661546;b=507325;opcode=000;
			#100	a=997827;b=-980246;opcode=010;
			#100	a=284549;b=219761;opcode=110;
			#100	a=442267;b=-344738;opcode=100;
			#100	a=604313;b=532818;opcode=010;
			#100	a=-23737;b=-285514;opcode=100;
			#100	a=-829973;b=-213710;opcode=111;
			#100	a=743213;b=100624;opcode=010;
			#100	a=804209;b=-259024;opcode=111;
			#100	a=-936331;b=748312;opcode=100;
			#100	a=501503;b=-729796;opcode=010;
			#100	a=875502;b=326702;opcode=100;
			#100	a=-197447;b=-95479;opcode=100;
			#100	a=913553;b=-480410;opcode=111;
			#100	a=-354896;b=-862741;opcode=001;
			#100	a=983622;b=-238232;opcode=111;
			#100	a=-170758;b=-408951;opcode=010;
			#100	a=-828021;b=-422595;opcode=010;
			#100	a=-380910;b=-635092;opcode=001;
			#100	a=31171;b=190097;opcode=000;
			#100	a=942776;b=768764;opcode=000;
			#100	a=429462;b=977845;opcode=001;
			#100	a=890929;b=169156;opcode=100;
			#100	a=-153809;b=135741;opcode=000;
			#100	a=-143561;b=-856828;opcode=001;
			#100	a=825371;b=756373;opcode=000;
			#100	a=-188303;b=-480481;opcode=000;
			#100	a=-544728;b=-923398;opcode=000;
			#100	a=-852049;b=-701337;opcode=010;
			#100	a=-745562;b=-180632;opcode=000;
			#100	a=-913544;b=-281907;opcode=010;
			#100	a=391408;b=-507422;opcode=010;
			#100	a=736843;b=537618;opcode=001;
			#100	a=-728587;b=-761810;opcode=001;
			#100	a=586967;b=44999;opcode=000;
			#100	a=205754;b=81223;opcode=001;
			#100	a=716523;b=-500059;opcode=010;
			#100	a=-818979;b=-527325;opcode=111;
			#100	a=-12213;b=272279;opcode=001;
			#100	a=-390463;b=-309149;opcode=001;
			#100	a=986388;b=381183;opcode=000;
			#100	a=-982384;b=-882304;opcode=100;
			#100	a=-158766;b=-811540;opcode=110;
			#100	a=146137;b=-760993;opcode=010;
			#100	a=750903;b=492983;opcode=110;
			#100	a=-317622;b=493300;opcode=001;
			#100	a=-262882;b=-874230;opcode=000;
			#100	a=-606921;b=566992;opcode=100;
			#100	a=184128;b=511362;opcode=000;
			#100	a=-757584;b=787613;opcode=100;
			#100	a=-5604;b=-242499;opcode=010;
			#100	a=-502229;b=-634141;opcode=010;
			#100	a=-435226;b=-561139;opcode=010;
			#100	a=387857;b=-272285;opcode=111;
			#100	a=-996700;b=757853;opcode=010;
			#100	a=770794;b=-237535;opcode=000;
			#100	a=-237258;b=-826340;opcode=110;
			#100	a=416077;b=343700;opcode=010;
			#100	a=17184;b=169666;opcode=110;
			#100	a=-60492;b=-196239;opcode=110;
			#100	a=-789244;b=504804;opcode=001;
			#100	a=-834716;b=-838060;opcode=100;
			#100	a=651100;b=-487186;opcode=001;
			#100	a=369843;b=666363;opcode=110;
			#100	a=-923675;b=228802;opcode=110;
			#100	a=910589;b=-464393;opcode=001;
			#100	a=581078;b=-948902;opcode=100;
			#100	a=-325580;b=514663;opcode=100;
			#100	a=-431206;b=888965;opcode=100;
			#100	a=496287;b=-419447;opcode=010;
			#100	a=-484566;b=-553136;opcode=010;
			#100	a=24930;b=-27553;opcode=110;
			#100	a=823016;b=-992964;opcode=010;
			#100	a=-145399;b=236577;opcode=001;
			#100	a=876227;b=369961;opcode=110;
			#100	a=-645209;b=-708921;opcode=110;
			#100	a=930001;b=-716836;opcode=100;
			#100	a=919228;b=-664104;opcode=001;
			#100	a=55232;b=361404;opcode=111;
			#100	a=537625;b=389715;opcode=001;
			#100	a=-307869;b=-256145;opcode=001;
			#100	a=837660;b=-959409;opcode=000;
			#100	a=63752;b=648125;opcode=110;
			#100	a=605291;b=296491;opcode=010;
			#100	a=-633212;b=-408491;opcode=100;
			#100	a=-302348;b=759376;opcode=010;
			#100	a=820382;b=473165;opcode=111;
			#100	a=687776;b=783802;opcode=100;
			#100	a=-144317;b=-640602;opcode=000;
			#100	a=804034;b=-766229;opcode=111;
			#100	a=-954494;b=-433982;opcode=110;
			#100	a=53001;b=176170;opcode=100;
			#100	a=-456343;b=556407;opcode=000;
			#100	a=-111181;b=696413;opcode=010;
			#100	a=-432381;b=167106;opcode=001;
			#100	a=839941;b=-184319;opcode=001;
			#100	a=555591;b=443760;opcode=100;
			#100	a=321956;b=-214467;opcode=010;
			#100	a=-930692;b=-468970;opcode=000;
			#100	a=-920196;b=-278667;opcode=001;
			#100	a=834877;b=-294342;opcode=001;
			#100	a=-150932;b=-412938;opcode=001;
			#100	a=540414;b=-906019;opcode=111;
			#100	a=-95872;b=624374;opcode=010;
			#100	a=-310360;b=-492689;opcode=111;
			#100	a=299791;b=171072;opcode=111;
			#100	a=-699568;b=-149285;opcode=000;
			#100	a=-403803;b=4567;opcode=100;
			#100	a=15155;b=358509;opcode=110;
			#100	a=-795829;b=708186;opcode=111;
			#100	a=656697;b=-778686;opcode=010;
			#100	a=318436;b=83732;opcode=111;
			#100	a=-760054;b=-886739;opcode=111;
			#100	a=-382819;b=-784585;opcode=110;
			#100	a=-421018;b=-241413;opcode=010;
			#100	a=-424509;b=448122;opcode=100;
			#100	a=-19672;b=738311;opcode=111;
			#100	a=-879846;b=917776;opcode=000;
			#100	a=657381;b=597141;opcode=000;
			#100	a=-665461;b=-634882;opcode=000;
			#100	a=589615;b=605795;opcode=111;
			#100	a=960713;b=819071;opcode=100;
			#100	a=-985515;b=-152252;opcode=100;
			#100	a=456715;b=787553;opcode=010;
			#100	a=-318300;b=387961;opcode=110;
			#100	a=456047;b=-542643;opcode=000;
			#100	a=266834;b=-689893;opcode=110;
			#100	a=-956727;b=-618915;opcode=110;
			#100	a=-277231;b=981722;opcode=001;
			#100	a=125757;b=652332;opcode=110;
			#100	a=-191499;b=446882;opcode=100;
			#100	a=449527;b=-46778;opcode=000;
			#100	a=789913;b=-527134;opcode=111;
			#100	a=-261977;b=77255;opcode=010;
			#100	a=46405;b=650608;opcode=111;
			#100	a=23931;b=127762;opcode=111;
			#100	a=772600;b=-569041;opcode=100;
			#100	a=200483;b=-112521;opcode=100;
			#100	a=-412497;b=900860;opcode=001;
			#100	a=646232;b=-681069;opcode=000;
			#100	a=-691037;b=2476;opcode=000;
			#100	a=837264;b=-259466;opcode=000;
			#100	a=-642098;b=515736;opcode=100;
			#100	a=676319;b=296487;opcode=000;
			#100	a=796620;b=113749;opcode=000;
			#100	a=-479536;b=221506;opcode=000;
			#100	a=29473;b=-111385;opcode=110;
			#100	a=-140809;b=573684;opcode=100;
			#100	a=-519146;b=352917;opcode=010;
			#100	a=825949;b=316419;opcode=001;
			#100	a=824801;b=788316;opcode=001;
			#100	a=-860070;b=-620381;opcode=000;
			#100	a=-403287;b=-115492;opcode=110;
			#100	a=518729;b=-429211;opcode=010;
			#100	a=-364053;b=-37404;opcode=110;
			#100	a=692639;b=-303840;opcode=010;
			#100	a=39481;b=-87816;opcode=110;
			#100	a=-234816;b=170819;opcode=111;
			#100	a=-391665;b=-360110;opcode=100;
			#100	a=-747917;b=-192326;opcode=111;
			#100	a=936635;b=491909;opcode=100;
			#100	a=-649764;b=-860672;opcode=110;
			#100	a=-421425;b=208345;opcode=010;
			#100	a=564634;b=-468049;opcode=000;
			#100	a=-598336;b=-644958;opcode=110;
			#100	a=235403;b=-245360;opcode=000;
			#100	a=226256;b=-928750;opcode=111;
			#100	a=66572;b=-558771;opcode=100;
			#100	a=-811186;b=-828099;opcode=111;
			#100	a=-315402;b=-958098;opcode=000;
			#100	a=-83666;b=-237680;opcode=100;
			#100	a=-512767;b=949753;opcode=100;
			#100	a=-842650;b=557450;opcode=111;
			#100	a=5425;b=-538887;opcode=110;
			#100	a=132076;b=-569871;opcode=110;
			#100	a=-133111;b=-334662;opcode=000;
			#100	a=349009;b=106762;opcode=110;
			#100	a=431116;b=-328291;opcode=111;
			#100	a=611330;b=655140;opcode=001;
			#100	a=541995;b=-452817;opcode=110;
			#100	a=-713259;b=315719;opcode=111;
			#100	a=-875070;b=894362;opcode=000;
			#100	a=446488;b=974552;opcode=000;
			#100	a=-296750;b=37303;opcode=111;
			#100	a=605378;b=734599;opcode=010;
			#100	a=107053;b=-300777;opcode=000;
			#100	a=291178;b=-395308;opcode=111;
			#100	a=660011;b=-484822;opcode=100;
			#100	a=-304907;b=127285;opcode=010;
			#100	a=280890;b=700409;opcode=110;
			#100	a=74085;b=-728762;opcode=000;
			#100	a=801384;b=644763;opcode=110;
			#100	a=-442476;b=-412762;opcode=010;
			#100	a=-230434;b=958472;opcode=010;
			#100	a=-201907;b=-885910;opcode=000;
			#100	a=576199;b=551723;opcode=000;
			#100	a=-683747;b=-197741;opcode=000;
			#100	a=376990;b=-987736;opcode=001;
			#100	a=-536622;b=-386509;opcode=000;
			#100	a=457550;b=-802650;opcode=010;
			#100	a=-288298;b=372451;opcode=111;
			#100	a=-251425;b=428221;opcode=010;
			#100	a=312286;b=91098;opcode=010;
			#100	a=-378628;b=-639197;opcode=001;
			#100	a=-548714;b=818704;opcode=001;
			#100	a=892811;b=-300253;opcode=111;
			#100	a=-298853;b=291391;opcode=010;
			#100	a=-274544;b=429051;opcode=111;
			#100	a=-344936;b=255162;opcode=010;
			#100	a=181256;b=421983;opcode=000;
			#100	a=421940;b=-678847;opcode=010;
			#100	a=-147217;b=-645629;opcode=111;
			#100	a=-483355;b=-315568;opcode=001;
			#100	a=-845110;b=-151424;opcode=010;
			#100	a=205396;b=-194474;opcode=110;
			#100	a=-574891;b=848145;opcode=001;
			#100	a=457129;b=72329;opcode=100;
			#100	a=-325326;b=-624017;opcode=001;
			#100	a=132461;b=638287;opcode=111;
			#100	a=309952;b=140007;opcode=110;
			#100	a=920274;b=-952847;opcode=001;
			#100	a=991966;b=-960144;opcode=111;
			#100	a=-861783;b=98752;opcode=001;
			#100	a=-340615;b=-275245;opcode=100;
			#100	a=-696673;b=-295342;opcode=001;
			#100	a=-460317;b=-76754;opcode=010;
			#100	a=874086;b=18306;opcode=000;
			#100	a=-708102;b=408976;opcode=111;
			#100	a=-278673;b=504229;opcode=100;
			#100	a=919085;b=-391108;opcode=010;
			#100	a=553196;b=294799;opcode=111;
			#100	a=829722;b=707646;opcode=111;
			#100	a=-181931;b=120364;opcode=001;
			#100	a=-838428;b=-444342;opcode=100;
			#100	a=-958518;b=403707;opcode=001;
			#100	a=-942084;b=53256;opcode=111;
			#100	a=-791566;b=462409;opcode=000;
			#100	a=-398641;b=419294;opcode=001;
			#100	a=771332;b=201175;opcode=100;
			#100	a=50101;b=55047;opcode=100;
			#100	a=-320223;b=-496413;opcode=111;
			#100	a=311352;b=-857926;opcode=000;
			#100	a=-837438;b=956388;opcode=010;
			#100	a=-912185;b=979281;opcode=111;
			#100	a=-613609;b=539705;opcode=110;
			#100	a=-411486;b=-434186;opcode=001;
			#100	a=-294056;b=-395984;opcode=110;
			#100	a=-118759;b=345549;opcode=111;
			#100	a=403698;b=-237476;opcode=100;
			#100	a=-302570;b=-627406;opcode=001;
			#100	a=542115;b=-652945;opcode=001;
			#100	a=-115947;b=874223;opcode=110;
			#100	a=211712;b=-479956;opcode=010;
			#100	a=750439;b=-794928;opcode=001;
			#100	a=-550529;b=-706546;opcode=100;
			#100	a=-625004;b=310823;opcode=010;
			#100	a=385460;b=-960576;opcode=001;
			#100	a=-140742;b=-702744;opcode=111;
			#100	a=834283;b=162627;opcode=010;
			#100	a=305329;b=-408432;opcode=001;
			#100	a=-46370;b=604804;opcode=100;
			#100	a=-410047;b=-294327;opcode=111;
			#100	a=-904516;b=-374568;opcode=100;
			#100	a=375150;b=84027;opcode=000;
			#100	a=904678;b=-221245;opcode=001;
			#100	a=-619042;b=789616;opcode=010;
			#100	a=-875975;b=-85469;opcode=010;
			#100	a=-966109;b=150805;opcode=110;
			#100	a=629869;b=36749;opcode=110;
			#100	a=-245575;b=291917;opcode=111;
			#100	a=142688;b=-490527;opcode=001;
			#100	a=-733538;b=986808;opcode=010;
			#100	a=-541680;b=-872917;opcode=000;
			#100	a=-866648;b=750542;opcode=111;
			#100	a=711993;b=-9832;opcode=100;
			#100	a=994219;b=-541401;opcode=111;
			#100	a=878289;b=-916513;opcode=111;
			#100	a=627092;b=479008;opcode=111;
			#100	a=-962410;b=-147281;opcode=000;
			#100	a=874525;b=945739;opcode=001;
			#100	a=-422811;b=-785839;opcode=111;
			#100	a=896842;b=208791;opcode=010;
			#100	a=-346754;b=-992238;opcode=100;
			#100	a=-805351;b=102791;opcode=111;
			#100	a=-335985;b=-684177;opcode=010;
			#100	a=606725;b=585944;opcode=100;
			#100	a=599627;b=875593;opcode=111;
			#100	a=486427;b=-435615;opcode=010;
			#100	a=-830313;b=-683354;opcode=111;
			#100	a=726396;b=697312;opcode=001;
			#100	a=267242;b=-467992;opcode=010;
			#100	a=-21303;b=526948;opcode=100;
			#100	a=-699340;b=495982;opcode=111;
			#100	a=515526;b=-710484;opcode=010;
			#100	a=923235;b=-550386;opcode=000;
			#100	a=-420492;b=702844;opcode=001;
			#100	a=-409765;b=-94077;opcode=010;
			#100	a=241315;b=775969;opcode=010;
			#100	a=-886657;b=85876;opcode=110;
			#100	a=-363751;b=-529706;opcode=111;
			#100	a=-37353;b=-928543;opcode=111;
			#100	a=505190;b=543019;opcode=010;
			#100	a=-305646;b=-815336;opcode=110;
			#100	a=52835;b=-30061;opcode=000;
			#100	a=23975;b=670823;opcode=010;
			#100	a=-968172;b=-228928;opcode=001;
			#100	a=-389582;b=157968;opcode=001;
			#100	a=-599434;b=216485;opcode=100;
			#100	a=-259753;b=317746;opcode=100;
			#100	a=-698435;b=194401;opcode=111;
			#100	a=-235096;b=-558687;opcode=100;
			#100	a=-464230;b=918151;opcode=000;
			#100	a=-855188;b=-638039;opcode=100;
			#100	a=-502435;b=243678;opcode=010;
			#100	a=895769;b=482622;opcode=000;
			#100	a=-421072;b=774007;opcode=010;
			#100	a=590807;b=487484;opcode=001;
			#100	a=145906;b=893258;opcode=110;
			#100	a=998341;b=-617777;opcode=100;
			#100	a=988964;b=-689314;opcode=100;
			#100	a=-962046;b=274082;opcode=000;
			#100	a=679622;b=-687505;opcode=100;
			#100	a=-547474;b=-390801;opcode=000;
			#100	a=-557457;b=-166556;opcode=110;
			#100	a=535857;b=-596656;opcode=100;
			#100	a=-655219;b=945832;opcode=110;
			#100	a=341216;b=53932;opcode=100;
			#100	a=-52232;b=497438;opcode=001;
			#100	a=478869;b=-619543;opcode=001;
			#100	a=-926465;b=563684;opcode=111;
			#100	a=978562;b=894474;opcode=111;
			#100	a=-532952;b=-830288;opcode=000;
			#100	a=140221;b=683027;opcode=000;
			#100	a=-250828;b=779559;opcode=100;
			#100	a=48114;b=-456565;opcode=001;
			#100	a=896483;b=157221;opcode=000;
			#100	a=399756;b=443512;opcode=010;
			#100	a=-283513;b=-799380;opcode=100;
			#100	a=-676500;b=997361;opcode=111;
			#100	a=975530;b=79642;opcode=001;
			#100	a=-560251;b=773248;opcode=010;
			#100	a=418653;b=584650;opcode=001;
			#100	a=756236;b=-338275;opcode=001;
			#100	a=-547959;b=-574727;opcode=010;
			#100	a=395760;b=694720;opcode=110;
			#100	a=-90589;b=-754714;opcode=111;
			#100	a=726081;b=95119;opcode=111;
			#100	a=-56026;b=-525242;opcode=001;
			#100	a=-963827;b=-466506;opcode=110;
			#100	a=955518;b=-609056;opcode=000;
			#100	a=684069;b=-535114;opcode=100;
			#100	a=329355;b=601939;opcode=110;
			#100	a=356921;b=-8280;opcode=010;
			#100	a=-725584;b=-294963;opcode=000;
			#100	a=742089;b=-381662;opcode=111;
			#100	a=211156;b=-381203;opcode=110;
			#100	a=-360317;b=958855;opcode=110;
			#100	a=175565;b=-719114;opcode=000;
			#100	a=9149;b=344913;opcode=110;
			#100	a=-141925;b=-283693;opcode=001;
			#100	a=-12992;b=-322153;opcode=110;
			#100	a=-988362;b=76036;opcode=001;
			#100	a=-703949;b=-902616;opcode=100;
			#100	a=-654414;b=214534;opcode=000;
			#100	a=-783261;b=-461405;opcode=100;
			#100	a=-397974;b=756562;opcode=010;
			#100	a=799746;b=-581606;opcode=111;
			#100	a=385816;b=252525;opcode=001;
			#100	a=-42760;b=641293;opcode=001;
			#100	a=-424296;b=774040;opcode=010;
			#100	a=713114;b=813406;opcode=000;
			#100	a=-839393;b=616191;opcode=001;
			#100	a=342650;b=-695933;opcode=000;
			#100	a=-742177;b=945027;opcode=110;
			#100	a=-82806;b=-448423;opcode=000;
			#100	a=-387639;b=-973112;opcode=110;
			#100	a=147057;b=-486747;opcode=100;
			#100	a=-526441;b=-521932;opcode=010;
			#100	a=-518069;b=-680758;opcode=100;
			#100	a=218451;b=396930;opcode=000;
			#100	a=-403944;b=93630;opcode=010;
			#100	a=692294;b=384877;opcode=110;
			#100	a=-626291;b=-39791;opcode=001;
			#100	a=599180;b=47855;opcode=100;
			#100	a=-249127;b=-425761;opcode=100;
			#100	a=451487;b=323674;opcode=110;
			#100	a=92419;b=31460;opcode=100;
			#100	a=-624616;b=486304;opcode=010;
			#100	a=147158;b=-35470;opcode=111;
			#100	a=676523;b=353850;opcode=110;
			#100	a=-614939;b=-163552;opcode=000;
			#100	a=-139502;b=753745;opcode=000;
			#100	a=-813721;b=-831686;opcode=110;
			#100	a=999177;b=-885140;opcode=100;
			#100	a=-876187;b=-999170;opcode=110;
			#100	a=770847;b=668930;opcode=001;
			#100	a=64614;b=-167471;opcode=110;
			#100	a=-416992;b=-363181;opcode=001;
			#100	a=162773;b=885734;opcode=100;
			#100	a=339128;b=-900242;opcode=001;
			#100	a=599465;b=71719;opcode=000;
			#100	a=-837395;b=25219;opcode=110;
			#100	a=-652349;b=-328735;opcode=010;
			#100	a=-728889;b=125089;opcode=000;
			#100	a=-918366;b=-227372;opcode=000;
			#100	a=-381375;b=754379;opcode=000;
			#100	a=194488;b=-766805;opcode=010;
			#100	a=-651976;b=-274562;opcode=100;
			#100	a=-319411;b=-461804;opcode=110;
			#100	a=-376473;b=470541;opcode=100;
			#100	a=-349541;b=554378;opcode=110;
			#100	a=107313;b=324360;opcode=110;
			#100	a=207788;b=411822;opcode=000;
			#100	a=989488;b=979992;opcode=000;
			#100	a=-667134;b=-62034;opcode=000;
			#100	a=342016;b=-56029;opcode=100;
			#100	a=861268;b=712175;opcode=000;
			#100	a=74543;b=209754;opcode=010;
			#100	a=-522719;b=396244;opcode=010;
			#100	a=-533028;b=984213;opcode=111;
			#100	a=-254840;b=308860;opcode=111;
			#100	a=214497;b=-400712;opcode=110;
			#100	a=-994818;b=-953173;opcode=110;
			#100	a=-775501;b=-768365;opcode=100;
			#100	a=-76132;b=726775;opcode=111;
			#100	a=-596979;b=-253062;opcode=111;
			#100	a=300471;b=-3778;opcode=010;
			#100	a=-739438;b=556314;opcode=000;
			#100	a=910395;b=-300693;opcode=000;
			#100	a=719362;b=-741075;opcode=110;
			#100	a=-954132;b=-697438;opcode=000;
			#100	a=-927140;b=935881;opcode=111;
			#100	a=245647;b=-226759;opcode=111;
			#100	a=935763;b=470331;opcode=000;
			#100	a=-306262;b=289824;opcode=010;
			#100	a=-287493;b=408684;opcode=110;
			#100	a=797307;b=821685;opcode=001;
			#100	a=-164515;b=-150048;opcode=010;
			#100	a=-232683;b=-588415;opcode=010;
			#100	a=-659259;b=230709;opcode=100;
			#100	a=653163;b=602142;opcode=100;
			#100	a=-742211;b=382768;opcode=010;
			#100	a=687688;b=414924;opcode=000;
			#100	a=433183;b=313660;opcode=010;
			#100	a=452917;b=984774;opcode=001;
			#100	a=858131;b=-416515;opcode=110;
			#100	a=-415236;b=152882;opcode=110;
			#100	a=-216363;b=-222369;opcode=100;
			#100	a=-886831;b=59901;opcode=001;
			#100	a=6913;b=-473604;opcode=100;
			#100	a=363794;b=29813;opcode=000;
			#100	a=354987;b=907654;opcode=001;
			#100	a=356734;b=-421334;opcode=001;
			#100	a=626268;b=-786696;opcode=000;
			#100	a=175814;b=-440451;opcode=010;
			#100	a=-595098;b=-37381;opcode=001;
			#100	a=500521;b=533869;opcode=000;
			#100	a=-962926;b=-151649;opcode=100;
			#100	a=-139909;b=839067;opcode=001;
			#100	a=102768;b=-486745;opcode=110;
			#100	a=-893513;b=692373;opcode=110;
			#100	a=373398;b=-674499;opcode=001;
			#100	a=92105;b=-671815;opcode=100;
			#100	a=-912;b=817595;opcode=010;
			#100	a=888042;b=373298;opcode=000;
			#100	a=-773540;b=-689404;opcode=110;
			#100	a=-741890;b=-83508;opcode=111;
			#100	a=-288598;b=-429674;opcode=000;
			#100	a=796926;b=-566144;opcode=110;
			#100	a=-736154;b=5447;opcode=110;
			#100	a=-762226;b=138164;opcode=001;
			#100	a=-771242;b=-338305;opcode=010;
			#100	a=175419;b=610871;opcode=100;
			#100	a=951498;b=915815;opcode=100;
			#100	a=482144;b=950137;opcode=110;
			#100	a=675627;b=99476;opcode=110;
			#100	a=-36012;b=831011;opcode=001;
			#100	a=-242943;b=-404759;opcode=010;
			#100	a=804167;b=167792;opcode=110;
			#100	a=-552714;b=249541;opcode=010;
			#100	a=-306991;b=-970036;opcode=010;
			#100	a=-634512;b=-618826;opcode=100;
			#100	a=-698718;b=-822004;opcode=100;
			#100	a=452432;b=-377163;opcode=000;
			#100	a=747743;b=363950;opcode=100;
			#100	a=44498;b=811565;opcode=111;
			#100	a=-358392;b=-323760;opcode=000;
			#100	a=-637064;b=-766928;opcode=100;
			#100	a=-508435;b=906720;opcode=100;
			#100	a=237267;b=514322;opcode=000;
			#100	a=-684226;b=-66034;opcode=111;
			#100	a=914089;b=-655399;opcode=001;
			#100	a=337409;b=-814908;opcode=010;
			#100	a=927060;b=-641554;opcode=000;
			#100	a=708851;b=-70949;opcode=000;
			#100	a=199052;b=289387;opcode=000;
			#100	a=882693;b=-709265;opcode=000;
			#100	a=-296027;b=-619345;opcode=001;
			#100	a=-359596;b=-926329;opcode=000;
			#100	a=484611;b=133552;opcode=000;
			#100	a=-580597;b=-167409;opcode=110;
			#100	a=113660;b=-911322;opcode=110;
			#100	a=217397;b=150025;opcode=000;
			#100	a=-357824;b=-157800;opcode=100;
			#100	a=-391963;b=-912146;opcode=010;
			#100	a=481482;b=-994694;opcode=110;
			#100	a=98009;b=-254012;opcode=001;
			#100	a=-991283;b=412499;opcode=000;
			#100	a=678301;b=-31891;opcode=000;
			#100	a=-285604;b=-408068;opcode=001;
			#100	a=-158798;b=138365;opcode=100;
			#100	a=-339027;b=476648;opcode=100;
			#100	a=-341890;b=-607907;opcode=000;
			#100	a=-901397;b=611841;opcode=010;
			#100	a=859311;b=-881513;opcode=010;
			#100	a=429298;b=-610728;opcode=010;
			#100	a=388630;b=-253056;opcode=111;
			#100	a=462259;b=702845;opcode=000;
			#100	a=-230378;b=398856;opcode=100;
			#100	a=53130;b=-94887;opcode=001;
			#100	a=79602;b=-62961;opcode=110;
			#100	a=-180206;b=-566978;opcode=000;
			#100	a=-896539;b=577358;opcode=000;
			#100	a=228742;b=137050;opcode=010;
			#100	a=483871;b=540420;opcode=001;
			#100	a=-426615;b=379624;opcode=110;
			#100	a=991844;b=-162677;opcode=110;
			#100	a=-717850;b=-771066;opcode=010;
			#100	a=461393;b=-102802;opcode=010;
			#100	a=24690;b=-275024;opcode=010;
			#100	a=-237762;b=272524;opcode=000;
			#100	a=39594;b=109173;opcode=100;
			#100	a=749815;b=-288420;opcode=000;
			#100	a=239592;b=481274;opcode=110;
			#100	a=-743189;b=-936497;opcode=010;
			#100	a=-427139;b=165198;opcode=001;
			#100	a=178284;b=431263;opcode=010;
			#100	a=-99755;b=-472809;opcode=110;
			#100	a=-471217;b=-463531;opcode=100;
			#100	a=-807533;b=-118051;opcode=111;
			#100	a=706106;b=-462967;opcode=010;
			#100	a=-916973;b=279197;opcode=010;
			#100	a=409465;b=-551682;opcode=001;
			#100	a=-142516;b=229787;opcode=110;
			#100	a=418729;b=-607271;opcode=110;
			#100	a=-847795;b=-982271;opcode=000;
			#100	a=309475;b=-100593;opcode=010;
			#100	a=-649031;b=519446;opcode=100;
			#100	a=-701178;b=-186619;opcode=100;
			#100	a=-486568;b=38895;opcode=010;
			#100	a=-860986;b=789385;opcode=001;
			#100	a=-15500;b=881667;opcode=000;
			#100	a=-84714;b=661808;opcode=111;
			#100	a=78931;b=495240;opcode=100;
			#100	a=-38972;b=-160818;opcode=100;
			#100	a=-924548;b=358184;opcode=111;
			#100	a=648957;b=735678;opcode=100;
			#100	a=812885;b=135830;opcode=000;
			#100	a=-968794;b=333201;opcode=111;
			#100	a=-612793;b=-93736;opcode=010;
			#100	a=-540981;b=-170806;opcode=100;
			#100	a=-225409;b=732741;opcode=110;
			#100	a=-242968;b=-38322;opcode=110;
			#100	a=327874;b=674388;opcode=100;
			#100	a=-649354;b=-283200;opcode=000;
			#100	a=-38197;b=-754;opcode=110;
			#100	a=99817;b=-451707;opcode=001;
			#100	a=-232091;b=755049;opcode=111;
			#100	a=-170558;b=839741;opcode=001;
			#100	a=-272256;b=485423;opcode=010;
			#100	a=252159;b=-233190;opcode=110;
			#100	a=843325;b=957523;opcode=110;
			#100	a=-305605;b=593394;opcode=010;
			#100	a=840529;b=185498;opcode=110;
			#100	a=498872;b=561003;opcode=000;
			#100	a=315346;b=356608;opcode=000;
			#100	a=137156;b=-416516;opcode=000;
			#100	a=290940;b=-317018;opcode=111;
			#100	a=-913565;b=794402;opcode=000;
			#100	a=665834;b=944833;opcode=010;
			#100	a=913957;b=-962289;opcode=110;
			#100	a=816670;b=73292;opcode=110;
			#100	a=-513924;b=-418863;opcode=100;
			#100	a=-944307;b=-412534;opcode=001;
			#100	a=15164;b=-141927;opcode=010;
			#100	a=781306;b=602591;opcode=001;
			#100	a=755144;b=-354518;opcode=111;
			#100	a=-145010;b=-981362;opcode=010;
			#100	a=461115;b=-761088;opcode=110;
			#100	a=80207;b=-427961;opcode=001;
			#100	a=683003;b=-778513;opcode=010;
			#100	a=-977046;b=37448;opcode=100;
			#100	a=177987;b=-743659;opcode=000;
			#100	a=-819765;b=963005;opcode=010;
			#100	a=-59030;b=292846;opcode=111;
			#100	a=-764058;b=260990;opcode=010;
			#100	a=46050;b=-889131;opcode=010;
			#100	a=-847805;b=717479;opcode=111;
			#100	a=351168;b=-356867;opcode=100;
			#100	a=660717;b=218900;opcode=001;
			#100	a=834584;b=-399647;opcode=111;
			#100	a=608748;b=953533;opcode=001;
			#100	a=-974651;b=-154731;opcode=010;
			#100	a=650044;b=682422;opcode=111;
			#100	a=548111;b=442202;opcode=010;
			#100	a=853726;b=560423;opcode=001;
			#100	a=234638;b=248621;opcode=111;
			#100	a=571879;b=532400;opcode=100;
			#100	a=191145;b=-684903;opcode=001;
			#100	a=-348226;b=658840;opcode=001;
			#100	a=815605;b=-529738;opcode=100;
			#100	a=-160272;b=964029;opcode=010;
			#100	a=-809673;b=-857324;opcode=001;
			#100	a=-450832;b=-182422;opcode=110;
			#100	a=-169194;b=8966;opcode=100;
			#100	a=-293115;b=-726348;opcode=001;
			#100	a=-607752;b=-938931;opcode=001;
			#100	a=-944309;b=-944024;opcode=100;
			#100	a=-12695;b=-584856;opcode=100;
			#100	a=449023;b=64571;opcode=000;
			#100	a=88872;b=102809;opcode=010;
			#100	a=223695;b=-808606;opcode=001;
			#100	a=191975;b=-872106;opcode=000;
			#100	a=-33674;b=-552845;opcode=111;
			#100	a=408429;b=-475923;opcode=000;
			#100	a=557468;b=250953;opcode=110;
			#100	a=946597;b=-897048;opcode=010;
			#100	a=-784640;b=361995;opcode=010;
			#100	a=48098;b=-128105;opcode=010;
			#100	a=128496;b=814999;opcode=110;
			#100	a=-177443;b=-597039;opcode=111;
			#100	a=596485;b=268772;opcode=000;
			#100	a=-884303;b=139354;opcode=000;
			#100	a=-94242;b=-316726;opcode=001;
			#100	a=-952966;b=878802;opcode=010;
			#100	a=-516725;b=-627202;opcode=110;
			#100	a=919725;b=-396905;opcode=000;
			#100	a=-366170;b=313256;opcode=010;
			#100	a=-502729;b=187498;opcode=001;
			#100	a=-56654;b=-109624;opcode=111;
			#100	a=945261;b=-636001;opcode=000;
			#100	a=-738894;b=677851;opcode=000;
			#100	a=-786658;b=-833075;opcode=000;
			#100	a=440453;b=-655200;opcode=000;
			#100	a=-186411;b=-936787;opcode=111;
			#100	a=944026;b=304166;opcode=010;
			#100	a=395066;b=-195778;opcode=001;
			#100	a=477127;b=-773016;opcode=000;
			#100	a=526850;b=-84689;opcode=001;
			#100	a=-132990;b=969447;opcode=110;
			#100	a=343770;b=526226;opcode=001;
			#100	a=-93303;b=192635;opcode=111;
			#100	a=563443;b=884162;opcode=110;
			#100	a=-537213;b=-771350;opcode=010;
			#100	a=967669;b=510765;opcode=100;
			#100	a=-223931;b=392681;opcode=111;
			#100	a=275036;b=743340;opcode=001;
			#100	a=-232531;b=-903264;opcode=001;
			#100	a=550437;b=17912;opcode=000;
			#100	a=393491;b=-173936;opcode=100;
			#100	a=43963;b=567730;opcode=001;
			#100	a=-226816;b=481875;opcode=010;
			#100	a=-646264;b=-488728;opcode=111;
			#100	a=-588155;b=997551;opcode=010;
			#100	a=897815;b=354795;opcode=110;
			#100	a=787638;b=942996;opcode=100;
			#100	a=814726;b=209410;opcode=111;
			#100	a=150750;b=-681041;opcode=110;
			#100	a=-745104;b=92317;opcode=001;
			#100	a=-153711;b=-484300;opcode=110;
			#100	a=-60955;b=-238526;opcode=000;
			#100	a=-285067;b=-312359;opcode=001;
			#100	a=71748;b=622684;opcode=010;
			#100	a=-823442;b=-137016;opcode=110;
			#100	a=-813461;b=-155652;opcode=111;
			#100	a=-221090;b=-166335;opcode=000;
			#100	a=-969021;b=862110;opcode=110;
			#100	a=-445697;b=-178378;opcode=100;
			#100	a=297971;b=323247;opcode=111;
			#100	a=-815442;b=-495397;opcode=100;
			#100	a=-845605;b=495822;opcode=010;
			#100	a=-609022;b=-921088;opcode=110;
			#100	a=-259760;b=-910931;opcode=000;
			#100	a=216738;b=-903022;opcode=110;
			#100	a=776078;b=96725;opcode=111;
			#100	a=-744351;b=-902569;opcode=001;
			#100	a=-379317;b=692230;opcode=110;
			#100	a=668697;b=-533770;opcode=110;
			#100	a=53876;b=239724;opcode=100;
			#100	a=149615;b=-438022;opcode=001;
			#100	a=504238;b=961431;opcode=001;
			#100	a=496036;b=326021;opcode=010;
			#100	a=182653;b=-462012;opcode=001;
			#100	a=426591;b=892202;opcode=001;
			#100	a=632004;b=-766390;opcode=001;
			#100	a=857581;b=418601;opcode=001;
			#100	a=346347;b=-585777;opcode=110;
			#100	a=-24848;b=-495155;opcode=111;
			#100	a=905354;b=871108;opcode=110;
			#100	a=-794518;b=816346;opcode=110;
			#100	a=599900;b=-694508;opcode=110;
			#100	a=-382837;b=-689390;opcode=010;
			#100	a=-375165;b=-573729;opcode=010;
			#100	a=-125884;b=66717;opcode=110;
			#100	a=-572497;b=-885577;opcode=111;
			#100	a=-437202;b=296183;opcode=001;
			#100	a=-730811;b=109977;opcode=001;
			#100	a=48237;b=-701447;opcode=001;
			#100	a=-934995;b=-967141;opcode=010;
			#100	a=-301737;b=554162;opcode=110;
			#100	a=566775;b=151749;opcode=000;
			#100	a=729948;b=163369;opcode=000;
			#100	a=712719;b=-477157;opcode=111;
			#100	a=762050;b=-19725;opcode=110;
			#100	a=195781;b=221585;opcode=110;
			#100	a=-118074;b=-397580;opcode=111;
			#100	a=-341231;b=271559;opcode=000;
			#100	a=197945;b=-571968;opcode=110;
			#100	a=-455349;b=849386;opcode=100;
			#100	a=-626280;b=-112602;opcode=000;
			#100	a=159091;b=-779120;opcode=010;
			#100	a=580049;b=497727;opcode=100;
			#100	a=-932415;b=-339933;opcode=110;
			#100	a=37141;b=-921834;opcode=010;
			#100	a=-611906;b=-901717;opcode=010;
			#100	a=671324;b=-683389;opcode=100;
			#100	a=-528766;b=957059;opcode=100;
			#100	a=-173073;b=100577;opcode=111;
			#100	a=-945515;b=-89042;opcode=110;
			#100	a=-275744;b=314471;opcode=001;
			#100	a=76750;b=360647;opcode=000;
			#100	a=-563180;b=-235685;opcode=111;
			#100	a=-410091;b=-671243;opcode=110;
			#100	a=-430079;b=-170597;opcode=110;
			#100	a=302587;b=904500;opcode=110;
			#100	a=8801;b=608305;opcode=000;
			#100	a=410543;b=-952943;opcode=000;
			#100	a=930268;b=-800951;opcode=110;
			#100	a=-771527;b=-39490;opcode=110;
			#100	a=448435;b=-863442;opcode=000;
			#100	a=277958;b=13318;opcode=100;
			#100	a=-417842;b=967146;opcode=010;
			#100	a=429665;b=-617362;opcode=100;
			#100	a=924036;b=213678;opcode=110;
			#100	a=-872534;b=216658;opcode=010;
			#100	a=-886850;b=-769902;opcode=001;
			#100	a=718231;b=-711007;opcode=000;
			#100	a=147698;b=-353163;opcode=000;
			#100	a=-683014;b=-317589;opcode=100;
			#100	a=-427593;b=567667;opcode=010;
			#100	a=205128;b=495002;opcode=100;
			#100	a=280580;b=-906862;opcode=100;
			#100	a=862597;b=-784476;opcode=010;
			#100	a=46850;b=496790;opcode=110;
			#100	a=151667;b=-902679;opcode=100;
			#100	a=603850;b=-666077;opcode=111;
			#100	a=73722;b=-803414;opcode=111;
			#100	a=-877978;b=384235;opcode=010;
			#100	a=745640;b=-422997;opcode=010;
			#100	a=183659;b=-547828;opcode=001;
			#100	a=-211017;b=450882;opcode=100;
			#100	a=857834;b=-102769;opcode=110;
			#100	a=20026;b=-577276;opcode=000;
			#100	a=876110;b=-850923;opcode=110;
			#100	a=-423657;b=-527653;opcode=110;
			#100	a=-5089;b=94485;opcode=111;
			#100	a=708;b=971654;opcode=110;
			#100	a=471886;b=287256;opcode=010;
			#100	a=154773;b=564125;opcode=110;
			#100	a=81060;b=-217085;opcode=001;
			#100	a=-263943;b=413000;opcode=111;
			#100	a=351903;b=-66027;opcode=010;
			#100	a=795066;b=-868063;opcode=100;
			#100	a=352414;b=-246261;opcode=010;
			#100	a=659008;b=-725492;opcode=001;
			#100	a=-695567;b=383200;opcode=110;
			#100	a=852393;b=-967842;opcode=010;
			#100	a=-854582;b=-166553;opcode=000;
			#100	a=-200839;b=-863751;opcode=001;
			#100	a=238860;b=507694;opcode=100;
			#100	a=-345734;b=637344;opcode=100;
			#100	a=-545312;b=-655153;opcode=111;
			#100	a=-689426;b=-547667;opcode=111;
			#100	a=-893916;b=723575;opcode=000;
			#100	a=92967;b=491378;opcode=100;
			#100	a=-696104;b=-679006;opcode=110;
			#100	a=166684;b=-325009;opcode=110;
			#100	a=614594;b=-491502;opcode=001;
			#100	a=-91473;b=-498995;opcode=110;
			#100	a=-908371;b=-544052;opcode=111;
			#100	a=285274;b=-842663;opcode=100;
			#100	a=659244;b=275796;opcode=001;
			#100	a=-744207;b=784445;opcode=001;
			#100	a=663272;b=-85224;opcode=100;
			#100	a=-923858;b=294416;opcode=010;
			#100	a=-195401;b=-637254;opcode=010;
			#100	a=380777;b=86152;opcode=001;
			#100	a=656331;b=268906;opcode=100;
			#100	a=-78355;b=-165950;opcode=110;
			#100	a=-572662;b=781173;opcode=010;
			#100	a=978648;b=-496900;opcode=001;
			#100	a=681998;b=-978244;opcode=010;
			#100	a=-143052;b=-39846;opcode=100;
			#100	a=-107757;b=-144437;opcode=010;
			#100	a=99100;b=-804736;opcode=000;
			#100	a=150902;b=-77713;opcode=000;
			#100	a=-536719;b=226732;opcode=010;
			#100	a=-45449;b=-936467;opcode=111;
			#100	a=-497570;b=-413592;opcode=000;
			#100	a=567163;b=-974566;opcode=001;
			#100	a=-93850;b=-964044;opcode=001;
			#100	a=-457734;b=160197;opcode=001;
			#100	a=-910694;b=-468992;opcode=000;
			#100	a=581595;b=611673;opcode=010;
			#100	a=84582;b=230408;opcode=001;
			#100	a=371173;b=-142754;opcode=000;
			#100	a=-987150;b=144552;opcode=111;
			#100	a=-49722;b=-114860;opcode=000;
			#100	a=-47105;b=-225730;opcode=000;
			#100	a=-895198;b=-333672;opcode=111;
			#100	a=772915;b=860187;opcode=111;
			#100	a=157193;b=-880624;opcode=000;
			#100	a=610517;b=203420;opcode=110;
			#100	a=302296;b=-37122;opcode=100;
			#100	a=-104808;b=-618603;opcode=100;
			#100	a=-262309;b=601583;opcode=000;
			#100	a=448338;b=81993;opcode=111;
			#100	a=-515365;b=-955513;opcode=111;
			#100	a=717637;b=-281763;opcode=000;
			#100	a=376194;b=966288;opcode=100;
			#100	a=497981;b=160838;opcode=001;
			#100	a=-753455;b=-532396;opcode=001;
			#100	a=-164871;b=-422002;opcode=001;
			#100	a=42834;b=181903;opcode=100;
			#100	a=-63055;b=470951;opcode=000;
			#100	a=-542330;b=-213398;opcode=001;
			#100	a=-375965;b=546424;opcode=001;
			#100	a=-846358;b=-713652;opcode=010;
			#100	a=-635748;b=826971;opcode=100;
			#100	a=621728;b=-702566;opcode=000;
			#100	a=-869776;b=26870;opcode=100;
			#100	a=55050;b=-150366;opcode=000;
			#100	a=213321;b=-943579;opcode=001;
			#100	a=-852757;b=-455960;opcode=111;
			#100	a=-952997;b=-70721;opcode=000;
			#100	a=138711;b=-128725;opcode=100;
			#100	a=-509441;b=-513824;opcode=001;
			#100	a=111440;b=-420807;opcode=001;
			#100	a=-174745;b=-611572;opcode=111;
			#100	a=760522;b=-924039;opcode=001;
			#100	a=540277;b=285814;opcode=001;
			#100	a=-146096;b=-297972;opcode=100;
			#100	a=-582511;b=-491745;opcode=000;
			#100	a=331777;b=-753786;opcode=010;
			#100	a=946864;b=-186213;opcode=110;
			#100	a=-253435;b=-292257;opcode=000;
			#100	a=-259811;b=-54167;opcode=001;
			#100	a=18575;b=-464928;opcode=111;
			#100	a=838894;b=43595;opcode=100;
			#100	a=621592;b=576565;opcode=111;
			#100	a=897917;b=7223;opcode=001;
			#100	a=-848632;b=58881;opcode=110;
			#100	a=-104093;b=537815;opcode=100;
			#100	a=-470544;b=705674;opcode=100;
			#100	a=101507;b=760854;opcode=111;
			#100	a=821809;b=648368;opcode=111;
			#100	a=481078;b=161249;opcode=110;
			#100	a=468186;b=835829;opcode=001;
			#100	a=745818;b=737844;opcode=110;
			#100	a=-443102;b=-323952;opcode=100;
			#100	a=738225;b=285211;opcode=110;
			#100	a=494069;b=875412;opcode=000;
			#100	a=-763784;b=851654;opcode=111;
			#100	a=-437512;b=-124905;opcode=111;
			#100	a=-790015;b=-969891;opcode=100;
			#100	a=94310;b=408367;opcode=010;
			#100	a=865025;b=-15984;opcode=100;
			#100	a=466500;b=-817462;opcode=000;
			#100	a=-314115;b=451616;opcode=010;
			#100	a=209155;b=689712;opcode=100;
			#100	a=-195887;b=296000;opcode=000;
			#100	a=-520087;b=-145651;opcode=000;
			#100	a=-494786;b=-344748;opcode=111;
			#100	a=-503975;b=-947439;opcode=010;
			#100	a=-215537;b=500459;opcode=111;
			#100	a=-886639;b=586340;opcode=001;
			#100	a=901764;b=210188;opcode=001;
			#100	a=875244;b=-870836;opcode=110;
			#100	a=958624;b=-878378;opcode=100;
			#100	a=60483;b=210148;opcode=001;
			#100	a=540068;b=324039;opcode=111;
			#100	a=-693222;b=642354;opcode=100;
			#100	a=-808923;b=-158300;opcode=001;
			#100	a=-105371;b=409096;opcode=010;
			#100	a=-31161;b=153192;opcode=100;
			#100	a=839159;b=-607267;opcode=010;
			#100	a=-271731;b=259374;opcode=110;
			#100	a=639302;b=-593803;opcode=000;
			#100	a=-870672;b=-296317;opcode=000;
			#100	a=-777046;b=-452392;opcode=000;
			#100	a=405874;b=-348049;opcode=000;
			#100	a=-370996;b=-792221;opcode=001;
			#100	a=-624757;b=827742;opcode=010;
			#100	a=-90777;b=-416888;opcode=001;
			#100	a=623016;b=-479055;opcode=001;
			#100	a=975704;b=-700520;opcode=100;
			#100	a=284570;b=-446155;opcode=000;
			#100	a=797601;b=706936;opcode=111;
			#100	a=-520362;b=-619837;opcode=100;
			#100	a=452629;b=616446;opcode=001;
			#100	a=652709;b=620728;opcode=111;
			#100	a=643633;b=482854;opcode=010;
			#100	a=-654036;b=711614;opcode=001;
			#100	a=176701;b=415222;opcode=100;
			#100	a=186966;b=437001;opcode=110;
			#100	a=363106;b=291131;opcode=111;
			#100	a=652914;b=202166;opcode=010;
			#100	a=-143450;b=68187;opcode=000;
			#100	a=536880;b=-787720;opcode=010;
			#100	a=834721;b=790512;opcode=111;
			#100	a=796517;b=-92707;opcode=111;
			#100	a=-484222;b=627149;opcode=100;
			#100	a=57795;b=681757;opcode=001;
			#100	a=-834104;b=-800848;opcode=111;
			#100	a=-949912;b=485856;opcode=110;
			#100	a=-409732;b=-420196;opcode=001;
			#100	a=441016;b=552829;opcode=100;
			#100	a=292638;b=-636965;opcode=000;
			#100	a=871883;b=701753;opcode=001;
			#100	a=183101;b=859638;opcode=000;
			#100	a=258500;b=688281;opcode=110;
			#100	a=666464;b=-302382;opcode=010;
			#100	a=-981103;b=-756497;opcode=001;
			#100	a=593660;b=948635;opcode=010;
			#100	a=702938;b=-59008;opcode=111;
			#100	a=244598;b=40509;opcode=100;
			#100	a=-862341;b=617528;opcode=001;
			#100	a=507807;b=-608623;opcode=000;
			#100	a=-211854;b=-512992;opcode=100;
			#100	a=55336;b=-62800;opcode=001;
			#100	a=-532068;b=-692066;opcode=001;
			#100	a=-450804;b=635405;opcode=000;
			#100	a=953460;b=152760;opcode=110;
			#100	a=858370;b=820953;opcode=001;
			#100	a=-76707;b=-336476;opcode=001;
			#100	a=-685024;b=773060;opcode=111;
			#100	a=-749186;b=959293;opcode=000;
			#100	a=-152557;b=436384;opcode=111;
			#100	a=-225840;b=-94912;opcode=100;
			#100	a=331397;b=-50267;opcode=001;
			#100	a=-887894;b=-665811;opcode=110;
			#100	a=873942;b=757362;opcode=001;
			#100	a=855070;b=72318;opcode=111;
			#100	a=71684;b=-96246;opcode=100;
			#100	a=627141;b=674409;opcode=001;
			#100	a=-519113;b=-561775;opcode=001;
			#100	a=135750;b=953609;opcode=010;
			#100	a=-3158;b=-279246;opcode=110;
			#100	a=208595;b=631300;opcode=010;
			#100	a=858675;b=-936961;opcode=110;
			#100	a=-313273;b=778490;opcode=000;
			#100	a=-468308;b=963731;opcode=100;
			#100	a=958402;b=820852;opcode=100;
			#100	a=369148;b=-457849;opcode=100;
			#100	a=-405338;b=-365081;opcode=111;
			#100	a=647758;b=966431;opcode=110;
			#100	a=80903;b=-276365;opcode=010;
			#100	a=791131;b=-497928;opcode=000;
			#100	a=-201320;b=462511;opcode=000;
			#100	a=144706;b=-529718;opcode=110;
			#100	a=-767594;b=-588885;opcode=000;
			#100	a=351496;b=-222804;opcode=110;
			#100	a=-353382;b=-96173;opcode=010;
			#100	a=-439583;b=-601804;opcode=010;
			#100	a=-875951;b=525733;opcode=110;
			#100	a=-951961;b=-9503;opcode=000;
			#100	a=468943;b=-480289;opcode=110;
			#100	a=-72620;b=554722;opcode=111;
			#100	a=319396;b=973948;opcode=000;
			#100	a=819170;b=420601;opcode=111;
			#100	a=-219464;b=335205;opcode=111;
			#100	a=727474;b=-307373;opcode=000;
			#100	a=901871;b=-550565;opcode=010;
			#100	a=510614;b=511531;opcode=001;
			#100	a=-271680;b=732738;opcode=111;
			#100	a=-218680;b=-820358;opcode=001;
			#100	a=504285;b=-867657;opcode=010;
			#100	a=204373;b=-124669;opcode=100;
			#100	a=-367977;b=-235046;opcode=010;
			#100	a=-749464;b=681726;opcode=100;
			#100	a=-444760;b=-748445;opcode=000;
			#100	a=350124;b=-580286;opcode=000;
			#100	a=28450;b=378209;opcode=110;
			#100	a=-848001;b=85601;opcode=010;
			#100	a=436329;b=-871414;opcode=110;
			#100	a=-10178;b=839657;opcode=010;
			#100	a=774588;b=-255096;opcode=001;
			#100	a=-428385;b=808575;opcode=001;
			#100	a=560810;b=-900052;opcode=111;
			#100	a=-38724;b=732082;opcode=100;
			#100	a=286666;b=441635;opcode=111;
			#100	a=90124;b=-655942;opcode=001;
			#100	a=85945;b=117591;opcode=000;
			#100	a=570658;b=-839798;opcode=110;
			#100	a=871774;b=247242;opcode=111;
			#100	a=-967556;b=-598901;opcode=111;
			#100	a=906861;b=-443433;opcode=100;
			#100	a=-918418;b=666857;opcode=010;
			#100	a=-779856;b=-202896;opcode=110;
			#100	a=364402;b=-432865;opcode=100;
			#100	a=-826333;b=476712;opcode=100;
			#100	a=-356717;b=950701;opcode=100;
			#100	a=215155;b=797477;opcode=100;
			#100	a=-907592;b=976912;opcode=100;
			#100	a=769730;b=714136;opcode=001;
			#100	a=-15225;b=-477784;opcode=000;
			#100	a=-962681;b=253593;opcode=001;
			#100	a=-155187;b=-359554;opcode=000;
			#100	a=892064;b=-924512;opcode=010;
			#100	a=-865025;b=-37332;opcode=001;
			#100	a=780699;b=-615696;opcode=111;
			#100	a=-842275;b=-278440;opcode=001;
			#100	a=151875;b=-36574;opcode=111;
			#100	a=-177002;b=-927890;opcode=001;
			#100	a=-602974;b=782887;opcode=111;
			#100	a=-772451;b=-139526;opcode=100;
			#100	a=-975144;b=-771691;opcode=110;
			#100	a=500709;b=372541;opcode=001;
			#100	a=-25844;b=113715;opcode=001;
			#100	a=31675;b=-115424;opcode=000;
			#100	a=-938827;b=-864890;opcode=110;
			#100	a=300394;b=583893;opcode=010;
			#100	a=305121;b=-593118;opcode=001;
			#100	a=-322676;b=591893;opcode=000;
			#100	a=328926;b=87247;opcode=100;
			#100	a=-384199;b=916170;opcode=100;
			#100	a=-72887;b=-809200;opcode=110;
			#100	a=-716953;b=-655624;opcode=110;
			#100	a=501325;b=513314;opcode=001;
			#100	a=-173563;b=-676983;opcode=111;
			#100	a=-490841;b=-989195;opcode=000;
			#100	a=259260;b=-364992;opcode=100;
			#100	a=-189092;b=37972;opcode=000;
			#100	a=-249346;b=431967;opcode=110;
			#100	a=280494;b=568411;opcode=111;
			#100	a=-71766;b=20847;opcode=000;
			#100	a=-47360;b=191123;opcode=111;
			#100	a=-434718;b=-555475;opcode=111;
			#100	a=-115718;b=-141709;opcode=100;
			#100	a=-23760;b=809320;opcode=001;
			#100	a=-720386;b=290140;opcode=110;
			#100	a=-164640;b=244612;opcode=110;
			#100	a=-154859;b=259611;opcode=111;
			#100	a=125695;b=63045;opcode=100;
			#100	a=865906;b=493038;opcode=010;
			#100	a=764511;b=12456;opcode=000;
			#100	a=-17038;b=-130952;opcode=111;
			#100	a=-962119;b=-949734;opcode=111;
			#100	a=-203639;b=691480;opcode=000;
			#100	a=761414;b=738208;opcode=001;
			#100	a=167802;b=61417;opcode=000;
			#100	a=-815753;b=185320;opcode=001;
			#100	a=780298;b=280039;opcode=111;
			#100	a=-777366;b=241161;opcode=001;
			#100	a=119267;b=-77494;opcode=000;
			#100	a=-487171;b=21795;opcode=000;
			#100	a=432271;b=-910799;opcode=111;
			#100	a=483487;b=328859;opcode=110;
			#100	a=-200968;b=-832183;opcode=110;
			#100	a=838464;b=-654181;opcode=111;
			#100	a=-760467;b=-944335;opcode=001;
			#100	a=698891;b=870292;opcode=001;
			#100	a=-965054;b=973333;opcode=010;
			#100	a=-664950;b=-942265;opcode=001;
			#100	a=-982843;b=455789;opcode=000;
			#100	a=-787779;b=624935;opcode=001;
			#100	a=876676;b=60297;opcode=100;
			#100	a=64532;b=942220;opcode=110;
			#100	a=736025;b=969421;opcode=100;
			#100	a=-622178;b=479857;opcode=100;
			#100	a=-651482;b=-196534;opcode=000;
			#100	a=-975107;b=-505710;opcode=100;
			#100	a=166522;b=624471;opcode=000;
			#100	a=746843;b=-232509;opcode=010;
			#100	a=-854674;b=745132;opcode=100;
			#100	a=12111;b=-877158;opcode=100;
			#100	a=291267;b=158470;opcode=000;
			#100	a=-957559;b=459070;opcode=110;
			#100	a=-825142;b=-747375;opcode=110;
			#100	a=652653;b=-739563;opcode=111;
			#100	a=-500742;b=-478034;opcode=100;
			#100	a=-302550;b=472806;opcode=001;
			#100	a=-913886;b=-850943;opcode=000;
			#100	a=615311;b=296977;opcode=000;
			#100	a=-592825;b=496693;opcode=100;
			#100	a=381005;b=-527794;opcode=111;
			#100	a=157200;b=118004;opcode=001;
			#100	a=-916396;b=-682297;opcode=100;
			#100	a=893109;b=285413;opcode=100;
			#100	a=198760;b=320800;opcode=001;
			#100	a=745766;b=640866;opcode=001;
			#100	a=-810690;b=187122;opcode=000;
			#100	a=245883;b=-461707;opcode=110;
			#100	a=-381155;b=-781951;opcode=100;
			#100	a=660366;b=-355475;opcode=110;
			#100	a=319838;b=-910085;opcode=001;
			#100	a=332900;b=73310;opcode=000;
			#100	a=750284;b=138965;opcode=010;
			#100	a=137567;b=806481;opcode=110;
			#100	a=-495530;b=908912;opcode=001;
			#100	a=-424049;b=799967;opcode=111;
			#100	a=607369;b=865869;opcode=010;
			#100	a=708446;b=902974;opcode=000;
			#100	a=551664;b=-189491;opcode=100;
			#100	a=730744;b=233392;opcode=111;
			#100	a=-268942;b=-161594;opcode=110;
			#100	a=-240361;b=-28524;opcode=100;
			#100	a=-887181;b=862614;opcode=000;
			#100	a=462358;b=458714;opcode=010;
			#100	a=-767453;b=818567;opcode=100;
			#100	a=200561;b=678919;opcode=110;
			#100	a=-153119;b=-408120;opcode=110;
			#100	a=-63730;b=-18683;opcode=001;
			#100	a=-41487;b=331870;opcode=110;
			#100	a=402667;b=685651;opcode=100;
			#100	a=736552;b=756928;opcode=110;
			#100	a=77722;b=277442;opcode=100;
			#100	a=874755;b=100884;opcode=100;
			#100	a=-792168;b=107466;opcode=000;
			#100	a=-129979;b=209839;opcode=111;
			#100	a=-401683;b=182530;opcode=010;
			#100	a=-795710;b=705879;opcode=000;
			#100	a=-567769;b=286974;opcode=111;
			#100	a=-987150;b=911483;opcode=110;
			#100	a=112591;b=74067;opcode=100;
			#100	a=885543;b=-970390;opcode=110;
			#100	a=-42789;b=449197;opcode=110;
			#100	a=271811;b=-878207;opcode=000;
			#100	a=751690;b=-411563;opcode=111;
			#100	a=-381867;b=-963761;opcode=111;
			#100	a=-590130;b=736469;opcode=100;
			#100	a=-677370;b=684711;opcode=111;
			#100	a=-370669;b=-134431;opcode=001;
			#100	a=-982409;b=-869135;opcode=010;
			#100	a=534772;b=-816566;opcode=000;
			#100	a=-891781;b=-538547;opcode=110;
			#100	a=-813611;b=-644228;opcode=000;
			#100	a=-983083;b=-298254;opcode=111;
			#100	a=-243315;b=-572576;opcode=001;
			#100	a=-991153;b=-9850;opcode=110;
			#100	a=-752278;b=-124460;opcode=000;
			#100	a=615401;b=931653;opcode=000;
			#100	a=863391;b=-135522;opcode=100;
			#100	a=-506357;b=-776503;opcode=000;
			#100	a=853524;b=-226703;opcode=100;
			#100	a=-754300;b=244376;opcode=010;
			#100	a=-586791;b=207019;opcode=001;
			#100	a=-954903;b=-221012;opcode=001;
			#100	a=872978;b=-798295;opcode=000;
			#100	a=359116;b=-981958;opcode=001;
			#100	a=-334366;b=922537;opcode=100;
			#100	a=404172;b=-806957;opcode=111;
			#100	a=-703997;b=-323107;opcode=000;
			#100	a=709746;b=-175166;opcode=001;
			#100	a=181107;b=-592249;opcode=000;
			#100	a=60501;b=-493532;opcode=110;
			#100	a=638028;b=486498;opcode=100;
			#100	a=-197617;b=104186;opcode=110;
			#100	a=318245;b=53501;opcode=000;
			#100	a=967205;b=-706403;opcode=110;
			#100	a=458374;b=-150106;opcode=000;
			#100	a=-134811;b=491667;opcode=000;
			#100	a=474601;b=110156;opcode=000;
			#100	a=-200126;b=-859959;opcode=111;
			#100	a=797192;b=-594146;opcode=111;
			#100	a=604961;b=342568;opcode=111;
			#100	a=-546534;b=523055;opcode=111;
			#100	a=623028;b=855974;opcode=001;
			#100	a=910132;b=-371386;opcode=111;
			#100	a=-306753;b=820029;opcode=111;
			#100	a=-89730;b=796421;opcode=100;
			#100	a=-311848;b=-629330;opcode=000;
			#100	a=739379;b=-530612;opcode=001;
			#100	a=-139367;b=588032;opcode=111;
			#100	a=80486;b=-578545;opcode=100;
			#100	a=-480953;b=-952052;opcode=000;
			#100	a=496309;b=-227273;opcode=010;
			#100	a=-310082;b=911799;opcode=000;
			#100	a=800970;b=-268089;opcode=111;
			#100	a=-988617;b=-183910;opcode=110;
			#100	a=307350;b=939251;opcode=100;
			#100	a=-115080;b=-225273;opcode=001;
			#100	a=122753;b=155847;opcode=111;
			#100	a=673462;b=41895;opcode=111;
			#100	a=764091;b=636031;opcode=001;
			#100	a=-142011;b=-429253;opcode=100;
			#100	a=-670811;b=-219392;opcode=100;
			#100	a=979701;b=721252;opcode=001;
			#100	a=-621188;b=609061;opcode=100;
			#100	a=482853;b=75172;opcode=001;
			#100	a=429365;b=418331;opcode=111;
			#100	a=210741;b=-533307;opcode=000;
			#100	a=-573038;b=360904;opcode=000;
			#100	a=-617888;b=-394635;opcode=110;
			#100	a=-583015;b=766906;opcode=010;
			#100	a=-154871;b=266293;opcode=110;
			#100	a=969076;b=-632249;opcode=111;
			#100	a=52947;b=211891;opcode=110;
			#100	a=-7841;b=718336;opcode=001;
			#100	a=37762;b=180803;opcode=010;
			#100	a=-267640;b=-881771;opcode=110;
			#100	a=-677759;b=-969412;opcode=010;
			#100	a=-124831;b=567814;opcode=111;
			#100	a=119417;b=220533;opcode=110;
			#100	a=-668309;b=-12191;opcode=100;
			#100	a=261888;b=348930;opcode=110;
			#100	a=873551;b=900053;opcode=110;
			#100	a=344248;b=696597;opcode=100;
			#100	a=-288474;b=-196784;opcode=111;
			#100	a=454304;b=955797;opcode=010;
			#100	a=-769595;b=584117;opcode=110;
			#100	a=661693;b=738016;opcode=000;
			#100	a=959316;b=730343;opcode=010;
			#100	a=387989;b=-350606;opcode=110;
			#100	a=-776522;b=-870035;opcode=100;
			#100	a=-158538;b=297200;opcode=010;
			#100	a=-72662;b=-625293;opcode=001;
			#100	a=572543;b=337784;opcode=001;
			#100	a=676130;b=-160044;opcode=110;
			#100	a=49155;b=-633869;opcode=100;
			#100	a=-184653;b=615277;opcode=110;
			#100	a=62168;b=-75505;opcode=111;
			#100	a=-572525;b=173835;opcode=001;
			#100	a=-906626;b=-611515;opcode=111;
			#100	a=-824167;b=26716;opcode=001;
			#100	a=935166;b=773494;opcode=000;
			#100	a=-390350;b=723238;opcode=100;
			#100	a=-177297;b=-677248;opcode=111;
			#100	a=-883013;b=-116645;opcode=100;
			#100	a=-353135;b=-962586;opcode=110;
			#100	a=-593367;b=928417;opcode=100;
			#100	a=-802400;b=886959;opcode=111;
			#100	a=415822;b=304990;opcode=110;
			#100	a=876881;b=-706474;opcode=000;
			#100	a=628676;b=852660;opcode=110;
			#100	a=-871753;b=323390;opcode=010;
			#100	a=904005;b=-437567;opcode=010;
			#100	a=-887133;b=209502;opcode=001;
			#100	a=-180102;b=191278;opcode=001;
			#100	a=-213821;b=-613364;opcode=110;
			#100	a=-18538;b=-401628;opcode=001;
			#100	a=-416776;b=395771;opcode=000;
			#100	a=145419;b=365243;opcode=010;
			#100	a=930847;b=359598;opcode=111;
			#100	a=352804;b=783863;opcode=111;
			#100	a=283971;b=-156035;opcode=001;
			#100	a=934870;b=-216545;opcode=001;
			#100	a=-946774;b=-982357;opcode=010;
			#100	a=-432177;b=804361;opcode=110;
			#100	a=-634467;b=-748210;opcode=100;
			#100	a=290057;b=433565;opcode=100;
			#100	a=695975;b=-390082;opcode=111;
			#100	a=-929291;b=-789775;opcode=111;
			#100	a=-89861;b=465855;opcode=001;
			#100	a=-542009;b=647810;opcode=100;
			#100	a=50172;b=-393842;opcode=010;
			#100	a=466445;b=433206;opcode=001;
			#100	a=173320;b=237319;opcode=110;
			#100	a=870480;b=472599;opcode=110;
			#100	a=-901908;b=-8104;opcode=001;
			#100	a=-858787;b=-680821;opcode=110;
			#100	a=-937762;b=576809;opcode=100;
			#100	a=647140;b=-864878;opcode=000;
			#100	a=106126;b=750776;opcode=010;
			#100	a=850418;b=623404;opcode=001;
			#100	a=184314;b=-515598;opcode=100;
			#100	a=-237958;b=-668552;opcode=100;
			#100	a=606553;b=-889813;opcode=001;
			#100	a=-474473;b=-122249;opcode=111;
			#100	a=-431406;b=-790927;opcode=001;
			#100	a=-243269;b=852012;opcode=111;
			#100	a=-969827;b=-866771;opcode=110;
			#100	a=545808;b=471828;opcode=001;
			#100	a=-4965;b=-726612;opcode=110;
			#100	a=-308910;b=165981;opcode=100;
			#100	a=905866;b=62898;opcode=110;
			#100	a=18816;b=-383176;opcode=110;
			#100	a=-79377;b=-717763;opcode=000;
			#100	a=573038;b=-894789;opcode=001;
			#100	a=-456324;b=-915179;opcode=000;
			#100	a=672975;b=887495;opcode=010;
			#100	a=595227;b=302564;opcode=000;
			#100	a=848694;b=-722648;opcode=100;
			#100	a=801485;b=-36537;opcode=111;
			#100	a=-566006;b=-180622;opcode=001;
			#100	a=915868;b=-366655;opcode=000;
			#100	a=843735;b=-156061;opcode=100;
			#100	a=881790;b=-829767;opcode=110;
			#100	a=-192194;b=-639308;opcode=100;
			#100	a=-176125;b=-580994;opcode=000;
			#100	a=-328090;b=498954;opcode=001;
			#100	a=416799;b=-734214;opcode=111;
			#100	a=449482;b=758663;opcode=001;
			#100	a=190477;b=-852749;opcode=010;
			#100	a=832403;b=724861;opcode=100;
			#100	a=-173392;b=51147;opcode=010;
			#100	a=750129;b=984385;opcode=001;
			#100	a=20549;b=-123960;opcode=010;
			#100	a=-863926;b=171097;opcode=001;
			#100	a=-562904;b=-622896;opcode=000;
			#100	a=-630992;b=516486;opcode=010;
			#100	a=118707;b=-303338;opcode=001;
			#100	a=68854;b=-689966;opcode=110;
			#100	a=515244;b=169298;opcode=001;
			#100	a=-150894;b=479442;opcode=110;
			#100	a=-297946;b=64692;opcode=000;
			#100	a=744967;b=-392115;opcode=001;
			#100	a=534759;b=-462329;opcode=001;
			#100	a=848730;b=832777;opcode=100;
			#100	a=274681;b=425645;opcode=100;
			#100	a=794153;b=-660425;opcode=001;
			#100	a=87696;b=949541;opcode=110;
			#100	a=-654148;b=-228277;opcode=010;
			#100	a=226807;b=-828543;opcode=100;
			#100	a=872247;b=743229;opcode=001;
			#100	a=980100;b=72914;opcode=100;
			#100	a=-458256;b=331732;opcode=110;
			#100	a=500633;b=134669;opcode=100;
			#100	a=-147459;b=888544;opcode=110;
			#100	a=-226822;b=472188;opcode=001;
			#100	a=711710;b=-491561;opcode=110;
			#100	a=922901;b=-85877;opcode=100;
			#100	a=-914457;b=-533504;opcode=001;
			#100	a=-27249;b=232866;opcode=000;
			#100	a=-463542;b=-513858;opcode=110;
			#100	a=767507;b=-229879;opcode=010;
			#100	a=148318;b=-196973;opcode=110;
			#100	a=1140;b=-33324;opcode=100;
			#100	a=-353534;b=739103;opcode=110;
			#100	a=532887;b=128068;opcode=010;
			#100	a=958018;b=-72211;opcode=010;
			#100	a=55586;b=913972;opcode=000;
			#100	a=195488;b=391252;opcode=111;
			#100	a=-877897;b=916415;opcode=111;
			#100	a=-45727;b=-942594;opcode=111;
			#100	a=858076;b=24587;opcode=110;
			#100	a=-672169;b=491304;opcode=001;
			#100	a=-817898;b=172269;opcode=100;
			#100	a=201068;b=-848902;opcode=010;
			#100	a=638454;b=873525;opcode=001;
			#100	a=-271808;b=-463959;opcode=100;
			#100	a=-312953;b=355993;opcode=111;
			#100	a=579299;b=683677;opcode=001;
			#100	a=717863;b=-14958;opcode=110;
			#100	a=588613;b=538159;opcode=110;
			#100	a=-399033;b=301728;opcode=110;
			#100	a=-383877;b=765996;opcode=111;
			#100	a=136536;b=107729;opcode=110;
			#100	a=87746;b=-97786;opcode=110;
			#100	a=586618;b=-674180;opcode=100;
			#100	a=-76826;b=902054;opcode=100;
			#100	a=-208196;b=-96264;opcode=001;
			#100	a=-990369;b=647456;opcode=010;
			#100	a=264055;b=800466;opcode=010;
			#100	a=-591532;b=845455;opcode=111;
			#100	a=-702284;b=673357;opcode=111;
			#100	a=-470198;b=927522;opcode=100;
			#100	a=-309439;b=41827;opcode=111;
			#100	a=962151;b=489573;opcode=010;
			#100	a=-422228;b=864056;opcode=110;
			#100	a=677524;b=817255;opcode=100;
			#100	a=-647861;b=-726317;opcode=000;
			#100	a=-285587;b=14157;opcode=001;
			#100	a=-930946;b=427950;opcode=100;
			#100	a=542357;b=438554;opcode=111;
			#100	a=200035;b=-486221;opcode=111;
			#100	a=693992;b=-620264;opcode=111;
			#100	a=40848;b=-553540;opcode=000;
			#100	a=659628;b=998246;opcode=000;
			#100	a=776420;b=145317;opcode=000;
			#100	a=445799;b=52873;opcode=111;
			#100	a=-209647;b=598831;opcode=000;
			#100	a=-201717;b=-142749;opcode=001;
			#100	a=363591;b=436018;opcode=100;
			#100	a=144716;b=-681459;opcode=000;
			#100	a=971899;b=-510081;opcode=110;
			#100	a=-358445;b=-702102;opcode=111;
			#100	a=686659;b=-35199;opcode=001;
			#100	a=-393344;b=-871946;opcode=110;
			#100	a=-879533;b=162138;opcode=001;
			#100	a=977965;b=-177730;opcode=001;
			#100	a=997426;b=-15366;opcode=110;
			#100	a=220446;b=975965;opcode=001;
			#100	a=178523;b=403717;opcode=100;
			#100	a=656062;b=-36984;opcode=111;
			#100	a=-908644;b=21918;opcode=111;
			#100	a=-839443;b=-915770;opcode=100;
			#100	a=-693008;b=-162931;opcode=110;
			#100	a=51642;b=-33931;opcode=100;
			#100	a=-956624;b=-756994;opcode=110;
			#100	a=869247;b=82515;opcode=110;
			#100	a=748593;b=-902523;opcode=010;
			#100	a=-779676;b=580480;opcode=111;
			#100	a=-758487;b=803657;opcode=000;
			#100	a=55075;b=-176669;opcode=000;
			#100	a=391691;b=582069;opcode=110;
			#100	a=95909;b=323824;opcode=100;
			#100	a=-811895;b=-312111;opcode=000;
			#100	a=-155876;b=525631;opcode=000;
			#100	a=173881;b=775776;opcode=010;
			#100	a=-338159;b=-160693;opcode=110;
			#100	a=601808;b=246627;opcode=110;
			#100	a=-655887;b=691710;opcode=000;
			#100	a=411630;b=-861986;opcode=010;
			#100	a=-201653;b=426;opcode=110;
			#100	a=-733026;b=859629;opcode=111;
			#100	a=40388;b=816651;opcode=001;
			#100	a=-318455;b=-129998;opcode=100;
			#100	a=-571771;b=922679;opcode=110;
			#100	a=-807695;b=996183;opcode=100;
			#100	a=-390187;b=227987;opcode=001;
			#100	a=396620;b=417933;opcode=100;
			#100	a=-660308;b=874784;opcode=010;
			#100	a=151992;b=521451;opcode=111;
			#100	a=-780507;b=-283027;opcode=110;
			#100	a=428549;b=-826778;opcode=001;
			#100	a=809801;b=-66252;opcode=010;
			#100	a=-992411;b=-531303;opcode=000;
			#100	a=-844251;b=-726060;opcode=010;
			#100	a=-645944;b=-152366;opcode=110;
			#100	a=722224;b=989492;opcode=100;
			#100	a=273086;b=396590;opcode=110;
			#100	a=136117;b=-161881;opcode=110;
			#100	a=-81580;b=245274;opcode=111;
			#100	a=-962501;b=-939635;opcode=111;
			#100	a=580471;b=378010;opcode=000;
			#100	a=-807745;b=828794;opcode=010;
			#100	a=200571;b=-649310;opcode=110;
			#100	a=17115;b=374420;opcode=001;
			#100	a=-508114;b=-99154;opcode=010;
			#100	a=-395590;b=665810;opcode=000;
			#100	a=-776611;b=593173;opcode=000;
			#100	a=-436357;b=-45944;opcode=010;
			#100	a=-712705;b=489893;opcode=000;
			#100	a=-632402;b=821323;opcode=010;
			#100	a=805544;b=-148646;opcode=001;
			#100	a=630668;b=-972769;opcode=100;
			#100	a=-722312;b=-831372;opcode=110;
			#100	a=-447318;b=875501;opcode=000;
			#100	a=980526;b=336948;opcode=110;
			#100	a=-499787;b=594203;opcode=010;
			#100	a=423734;b=-360548;opcode=001;
			#100	a=-881996;b=-893818;opcode=001;
			#100	a=-80822;b=423951;opcode=110;
			#100	a=794880;b=338836;opcode=111;
			#100	a=574560;b=561947;opcode=001;
			#100	a=-68999;b=-850793;opcode=111;
			#100	a=-279336;b=-40271;opcode=110;
			#100	a=741160;b=112274;opcode=100;
			#100	a=422753;b=-1271;opcode=001;
			#100	a=-766779;b=84774;opcode=000;
			#100	a=885345;b=-910588;opcode=001;
			#100	a=463921;b=-725621;opcode=110;
			#100	a=345754;b=565568;opcode=100;
			#100	a=597143;b=945021;opcode=110;
			#100	a=-133086;b=-383788;opcode=010;
			#100	a=913104;b=-398839;opcode=010;
			#100	a=276838;b=139973;opcode=111;
			#100	a=428885;b=942610;opcode=100;
			#100	a=747656;b=133780;opcode=000;
			#100	a=905812;b=-524543;opcode=001;
			#100	a=686283;b=563572;opcode=000;
			#100	a=-430611;b=87718;opcode=110;
			#100	a=-33076;b=273780;opcode=001;
			#100	a=-473177;b=369513;opcode=100;
			#100	a=-320241;b=-174178;opcode=000;
			#100	a=217750;b=-421459;opcode=000;
			#100	a=-958489;b=-735062;opcode=001;
			#100	a=173990;b=-680338;opcode=010;
			#100	a=483442;b=610323;opcode=010;
			#100	a=-291592;b=449655;opcode=000;
			#100	a=147897;b=349969;opcode=110;
			#100	a=815228;b=-603245;opcode=100;
			#100	a=89792;b=863703;opcode=100;
			#100	a=646287;b=-132169;opcode=100;
			#100	a=-97461;b=231662;opcode=100;
			#100	a=-954095;b=432323;opcode=111;
			#100	a=-632077;b=698922;opcode=100;
			#100	a=-722336;b=555941;opcode=110;
			#100	a=682980;b=-496084;opcode=111;
			#100	a=-350595;b=542083;opcode=111;
			#100	a=-328656;b=140514;opcode=001;
			#100	a=351821;b=600521;opcode=100;
			#100	a=376307;b=265548;opcode=110;
			#100	a=-512515;b=-48434;opcode=010;
			#100	a=-546331;b=577274;opcode=000;
			#100	a=536629;b=-20351;opcode=111;
			#100	a=-806317;b=245666;opcode=100;
			#100	a=-4561;b=-913690;opcode=111;
			#100	a=99538;b=873987;opcode=110;
			#100	a=938339;b=388143;opcode=110;
			#100	a=7373;b=-850156;opcode=100;
			#100	a=751929;b=306165;opcode=001;
			#100	a=-729407;b=-500268;opcode=100;
			#100	a=912163;b=-812920;opcode=111;
			#100	a=37433;b=-848633;opcode=001;
			#100	a=825031;b=-832767;opcode=000;
			#100	a=666669;b=496357;opcode=001;
			#100	a=343477;b=791255;opcode=000;
			#100	a=-328071;b=-99187;opcode=111;
			#100	a=-833604;b=217313;opcode=111;
			#100	a=-932874;b=-421345;opcode=110;
			#100	a=489881;b=872498;opcode=111;
			#100	a=-196720;b=-50671;opcode=111;
			#100	a=904711;b=-314791;opcode=100;
			#100	a=398219;b=-861667;opcode=000;
			#100	a=-930380;b=-495510;opcode=010;
			#100	a=736050;b=-221604;opcode=110;
			#100	a=862264;b=-42094;opcode=000;
			#100	a=-541179;b=-905445;opcode=111;
			#100	a=-661230;b=-50049;opcode=001;
			#100	a=-88864;b=-115241;opcode=010;
			#100	a=804731;b=-313195;opcode=111;
			#100	a=-36091;b=243006;opcode=110;
			#100	a=427396;b=-139947;opcode=001;
			#100	a=-555188;b=-110936;opcode=111;
			#100	a=-389148;b=326517;opcode=010;
			#100	a=-392924;b=670167;opcode=010;
			#100	a=994525;b=-650693;opcode=111;
			#100	a=-432248;b=924549;opcode=110;
			#100	a=-701460;b=-775611;opcode=000;
			#100	a=-592329;b=966778;opcode=111;
			#100	a=-937502;b=84019;opcode=000;
			#100	a=720232;b=874402;opcode=010;
			#100	a=-645119;b=-220257;opcode=010;
			#100	a=236970;b=486163;opcode=100;
			#100	a=-472842;b=-262511;opcode=110;
			#100	a=985756;b=632887;opcode=110;
			#100	a=-934240;b=-679865;opcode=010;
			#100	a=506165;b=866354;opcode=000;
			#100	a=-680394;b=80462;opcode=001;
			#100	a=195710;b=-308988;opcode=111;
			#100	a=139216;b=616406;opcode=110;
			#100	a=-395048;b=620458;opcode=000;
			#100	a=920252;b=163502;opcode=000;
			#100	a=765044;b=-184093;opcode=111;
			#100	a=-376085;b=-546086;opcode=110;
			#100	a=699466;b=215614;opcode=010;
			#100	a=525066;b=-725559;opcode=010;
			#100	a=-962047;b=-109418;opcode=111;
			#100	a=-560985;b=-115520;opcode=001;
			#100	a=130596;b=853620;opcode=000;
			#100	a=186465;b=-832578;opcode=100;
			#100	a=-339394;b=802060;opcode=100;
			#100	a=-16099;b=-337845;opcode=001;
			#100	a=-857123;b=979266;opcode=100;
			#100	a=-370447;b=644579;opcode=010;
			#100	a=44171;b=949933;opcode=100;
			#100	a=648523;b=-406501;opcode=110;
			#100	a=567246;b=-6636;opcode=001;
			#100	a=-696826;b=-8309;opcode=111;
			#100	a=-521872;b=320673;opcode=100;
			#100	a=-423524;b=194736;opcode=100;
			#100	a=800325;b=675437;opcode=100;
			#100	a=115493;b=559813;opcode=111;
			#100	a=331832;b=-776411;opcode=111;
			#100	a=-42542;b=-927773;opcode=100;
			#100	a=916045;b=697928;opcode=100;
			#100	a=-422768;b=227230;opcode=000;
			#100	a=-888129;b=883658;opcode=110;
			#100	a=-140493;b=-890399;opcode=010;
			#100	a=145953;b=-520764;opcode=001;
			#100	a=-914161;b=-298672;opcode=111;
			#100	a=960899;b=-739167;opcode=110;
			#100	a=-372012;b=-790884;opcode=001;
			#100	a=165213;b=223604;opcode=010;
			#100	a=981550;b=509311;opcode=111;
			#100	a=471174;b=996833;opcode=010;
			#100	a=647608;b=711894;opcode=111;
			#100	a=679222;b=-827703;opcode=001;
			#100	a=-931511;b=640307;opcode=000;
			#100	a=-768552;b=716716;opcode=001;
			#100	a=-60087;b=909189;opcode=111;
			#100	a=-51286;b=564929;opcode=110;
			#100	a=-838871;b=-230586;opcode=000;
			#100	a=391243;b=-90949;opcode=001;
			#100	a=948341;b=713425;opcode=111;
			#100	a=180683;b=-878181;opcode=000;
			#100	a=290889;b=-247130;opcode=110;
			#100	a=-348050;b=836983;opcode=001;
			#100	a=880930;b=507196;opcode=100;
			#100	a=-191042;b=-924160;opcode=110;
			#100	a=-482091;b=-125279;opcode=001;
			#100	a=389226;b=781028;opcode=100;
			#100	a=-781057;b=550434;opcode=100;
			#100	a=-79254;b=48091;opcode=100;
			#100	a=955980;b=571824;opcode=001;
			#100	a=46822;b=-393598;opcode=111;
			#100	a=-639;b=374568;opcode=111;
			#100	a=-187440;b=-803145;opcode=100;
			#100	a=92815;b=-940464;opcode=010;
			#100	a=695338;b=-408731;opcode=110;
			#100	a=439011;b=-293695;opcode=110;
			#100	a=-134165;b=11136;opcode=000;
			#100	a=484878;b=292447;opcode=110;
			#100	a=391857;b=-766538;opcode=110;
			#100	a=-172750;b=799269;opcode=111;
			#100	a=933075;b=-125700;opcode=001;
			#100	a=-236635;b=221188;opcode=000;
			#100	a=28953;b=-322137;opcode=100;
			#100	a=835611;b=-542273;opcode=111;
			#100	a=312984;b=-595898;opcode=010;
			#100	a=173180;b=127171;opcode=111;
			#100	a=145885;b=61989;opcode=010;
			#100	a=-739290;b=-404371;opcode=111;
			#100	a=-708224;b=-738793;opcode=110;
			#100	a=738395;b=264763;opcode=001;
			#100	a=-535663;b=357297;opcode=001;
			#100	a=-639870;b=-14099;opcode=110;
			#100	a=-811069;b=-960543;opcode=111;
			#100	a=-251445;b=-41384;opcode=100;
			#100	a=903140;b=475594;opcode=100;
			#100	a=606391;b=-519468;opcode=110;
			#100	a=27166;b=-108229;opcode=110;
			#100	a=-856789;b=302621;opcode=000;
			#100	a=572979;b=823106;opcode=000;
			#100	a=-394777;b=678012;opcode=111;
			#100	a=-566034;b=-486345;opcode=000;
			#100	a=945109;b=-78332;opcode=000;
			#100	a=-78492;b=-863799;opcode=100;
			#100	a=383355;b=-861799;opcode=000;
			#100	a=194037;b=381440;opcode=110;
			#100	a=-46155;b=-599862;opcode=001;
			#100	a=357030;b=115677;opcode=010;
			#100	a=970160;b=-627430;opcode=111;
			#100	a=-787251;b=-211725;opcode=100;
			#100	a=-41400;b=-767393;opcode=100;
			#100	a=580957;b=-672960;opcode=111;
			#100	a=510983;b=754234;opcode=000;
			#100	a=-279667;b=533704;opcode=010;
			#100	a=748300;b=-118819;opcode=010;
			#100	a=-646926;b=-644134;opcode=111;
			#100	a=-526779;b=-412655;opcode=001;
			#100	a=32174;b=-650721;opcode=001;
			#100	a=-863306;b=-468833;opcode=000;
			#100	a=914466;b=999351;opcode=100;
			#100	a=729189;b=-47050;opcode=001;
			#100	a=-922595;b=-965549;opcode=100;
			#100	a=-462146;b=-140333;opcode=010;
			#100	a=783380;b=634979;opcode=100;
			#100	a=-942369;b=-408876;opcode=010;
			#100	a=504707;b=393724;opcode=010;
			#100	a=-106074;b=-184250;opcode=010;
			#100	a=936430;b=-705933;opcode=010;
			#100	a=375048;b=130467;opcode=110;
			#100	a=916131;b=-229365;opcode=100;
			#100	a=861842;b=349725;opcode=010;
			#100	a=948243;b=130255;opcode=111;
			#100	a=-246618;b=-127620;opcode=010;
			#100	a=167602;b=64904;opcode=110;
			#100	a=919635;b=827695;opcode=100;
			#100	a=434772;b=-151174;opcode=100;
			#100	a=777232;b=814976;opcode=001;
			#100	a=985229;b=955463;opcode=001;
			#100	a=-61323;b=-658829;opcode=110;
			#100	a=66202;b=906600;opcode=010;
			#100	a=875977;b=-86898;opcode=001;
			#100	a=911790;b=-673160;opcode=000;
			#100	a=131054;b=-416119;opcode=001;
			#100	a=238672;b=-403993;opcode=110;
			#100	a=-865073;b=485892;opcode=001;
			#100	a=-821812;b=974294;opcode=110;
			#100	a=734445;b=997197;opcode=010;
			#100	a=647831;b=797048;opcode=100;
			#100	a=204757;b=-64307;opcode=111;
			#100	a=-127324;b=626083;opcode=001;
			#100	a=746707;b=-661028;opcode=001;
			#100	a=-245413;b=-797846;opcode=000;
			#100	a=-376061;b=-922736;opcode=110;
			#100	a=-203916;b=416494;opcode=111;
			#100	a=-7323;b=-544561;opcode=100;
			#100	a=105282;b=-363920;opcode=010;
			#100	a=-853592;b=413557;opcode=000;
			#100	a=449905;b=-471908;opcode=000;
			#100	a=825210;b=-852930;opcode=010;
			#100	a=-102979;b=783334;opcode=000;
			#100	a=-428593;b=656734;opcode=100;
			#100	a=-78501;b=15449;opcode=100;
			#100	a=-995285;b=-244468;opcode=100;
			#100	a=-457450;b=-436338;opcode=010;
			#100	a=569407;b=175927;opcode=100;
			#100	a=654880;b=149445;opcode=001;
			#100	a=-467998;b=739916;opcode=000;
			#100	a=373715;b=-68066;opcode=111;
			#100	a=-588325;b=-693340;opcode=000;
			#100	a=-733188;b=623366;opcode=111;
			#100	a=-864885;b=299545;opcode=100;
			#100	a=802560;b=550816;opcode=010;
			#100	a=198712;b=-648278;opcode=010;
			#100	a=-38252;b=860695;opcode=100;
			#100	a=423591;b=-242741;opcode=000;
			#100	a=-623311;b=-143820;opcode=111;
			#100	a=819425;b=365621;opcode=110;
			#100	a=594880;b=935930;opcode=110;
			#100	a=-22595;b=673962;opcode=000;
			#100	a=325842;b=-579556;opcode=100;
			#100	a=-197560;b=550489;opcode=110;
			#100	a=-992773;b=-786200;opcode=100;
			#100	a=-39526;b=128118;opcode=100;
			#100	a=-40852;b=917744;opcode=000;
			#100	a=487411;b=387910;opcode=010;
			#100	a=-52617;b=391735;opcode=010;
			#100	a=87941;b=975152;opcode=111;
			#100	a=-701886;b=-21516;opcode=110;
			#100	a=-43021;b=851067;opcode=010;
			#100	a=-816005;b=-560618;opcode=001;
			#100	a=890299;b=-727441;opcode=000;
			#100	a=958598;b=-383414;opcode=001;
			#100	a=849661;b=-432372;opcode=010;
			#100	a=120698;b=-230418;opcode=110;
			#100	a=138166;b=619411;opcode=000;
			#100	a=83968;b=-513032;opcode=001;
			#100	a=-860064;b=404765;opcode=111;
			#100	a=-602255;b=-386813;opcode=110;
			#100	a=293545;b=-288128;opcode=111;
			#100	a=346031;b=304185;opcode=111;
			#100	a=-308066;b=747392;opcode=010;
			#100	a=-520532;b=56427;opcode=111;
			#100	a=554031;b=-632447;opcode=111;
			#100	a=808155;b=-846199;opcode=000;
			#100	a=-900075;b=-346885;opcode=100;
			#100	a=-541395;b=-33051;opcode=110;
			#100	a=93720;b=-669733;opcode=110;
			#100	a=-595186;b=-348878;opcode=111;
			#100	a=-811686;b=-165203;opcode=000;
			#100	a=126949;b=399329;opcode=001;
			#100	a=947568;b=-540584;opcode=100;
			#100	a=-90631;b=886540;opcode=100;
			#100	a=994769;b=193548;opcode=111;
			#100	a=-214386;b=823233;opcode=100;
			#100	a=-218104;b=-147177;opcode=000;
			#100	a=-421456;b=-516077;opcode=000;
			#100	a=-602543;b=-328415;opcode=100;
			#100	a=173704;b=-544965;opcode=100;
			#100	a=-663500;b=-356496;opcode=100;
			#100	a=-337329;b=-49489;opcode=010;
			#100	a=-829299;b=-132292;opcode=110;
			#100	a=99685;b=976748;opcode=100;
			#100	a=-806458;b=-782064;opcode=001;
			#100	a=209935;b=113107;opcode=111;
			#100	a=-753309;b=12694;opcode=001;
			#100	a=786517;b=-321155;opcode=100;
			#100	a=5781;b=73026;opcode=010;
			#100	a=-601423;b=551669;opcode=001;
			#100	a=-94537;b=249539;opcode=000;
			#100	a=196095;b=152442;opcode=111;
			#100	a=-789089;b=-756213;opcode=010;
			#100	a=41756;b=-834536;opcode=000;
			#100	a=448335;b=431461;opcode=001;
			#100	a=466450;b=148464;opcode=001;
			#100	a=-780094;b=81098;opcode=000;
			#100	a=273436;b=319330;opcode=000;
			#100	a=578774;b=710134;opcode=000;
			#100	a=664222;b=481937;opcode=100;
			#100	a=122086;b=-378066;opcode=010;
			#100	a=-565970;b=63137;opcode=001;
			#100	a=-138913;b=356675;opcode=010;
			#100	a=-326589;b=300969;opcode=010;
			#100	a=258452;b=43178;opcode=111;
			#100	a=-403135;b=34461;opcode=100;
			#100	a=-360179;b=302905;opcode=100;
			#100	a=-523320;b=811223;opcode=100;
			#100	a=-429311;b=2600;opcode=111;
			#100	a=-189118;b=-748381;opcode=010;
			#100	a=-777944;b=-824915;opcode=001;
			#100	a=919864;b=361172;opcode=111;
			#100	a=-640862;b=-165908;opcode=100;
			#100	a=-896363;b=-299348;opcode=100;
			#100	a=-761427;b=478843;opcode=010;
			#100	a=-129690;b=107008;opcode=110;
			#100	a=994009;b=710663;opcode=000;
			#100	a=944260;b=336887;opcode=111;
			#100	a=142340;b=60791;opcode=010;
			#100	a=-684998;b=-470881;opcode=110;
			#100	a=-207853;b=573171;opcode=100;
			#100	a=-97656;b=140229;opcode=100;
			#100	a=342677;b=-524744;opcode=100;
			#100	a=-248873;b=-806515;opcode=010;
			#100	a=-961684;b=-326605;opcode=000;
			#100	a=-853512;b=-332389;opcode=000;
			#100	a=884250;b=-969371;opcode=110;
			#100	a=-409581;b=-954622;opcode=110;
			#100	a=129448;b=-234675;opcode=111;
			#100	a=-912370;b=-571186;opcode=001;
			#100	a=1825;b=141566;opcode=100;
			#100	a=-421994;b=-843920;opcode=100;
			#100	a=384880;b=99770;opcode=111;
			#100	a=-280191;b=-969318;opcode=000;
			#100	a=324718;b=962439;opcode=001;
			#100	a=-838799;b=-36920;opcode=111;
			#100	a=755454;b=647006;opcode=100;
			#100	a=493629;b=516142;opcode=110;
			#100	a=-801695;b=-961452;opcode=111;
			#100	a=-209335;b=680677;opcode=010;
			#100	a=-868246;b=-922247;opcode=110;
			#100	a=979318;b=487281;opcode=110;
			#100	a=-398469;b=-366010;opcode=110;
			#100	a=-716233;b=725438;opcode=111;
			#100	a=-581473;b=-467486;opcode=100;
			#100	a=129574;b=-739013;opcode=100;
			#100	a=49876;b=-930546;opcode=000;
			#100	a=-63533;b=144093;opcode=110;
			#100	a=872840;b=-223398;opcode=110;
			#100	a=787017;b=472084;opcode=001;
			#100	a=854438;b=-926468;opcode=010;
			#100	a=642172;b=703047;opcode=100;
			#100	a=493166;b=152497;opcode=111;
			#100	a=447044;b=894562;opcode=001;
			#100	a=-542149;b=275899;opcode=001;
			#100	a=223062;b=268464;opcode=010;
			#100	a=11687;b=586256;opcode=010;
			#100	a=44455;b=-362213;opcode=010;
			#100	a=960466;b=568388;opcode=110;
			#100	a=-724344;b=-670433;opcode=010;
			#100	a=-665439;b=-703352;opcode=001;
			#100	a=-717938;b=832615;opcode=110;
			#100	a=365157;b=403998;opcode=000;
			#100	a=983070;b=-478323;opcode=100;
			#100	a=76348;b=114637;opcode=000;
			#100	a=67148;b=544351;opcode=001;
			#100	a=-950630;b=-234182;opcode=100;
			#100	a=-145355;b=-622179;opcode=010;
			#100	a=951593;b=-672525;opcode=001;
			#100	a=745528;b=866611;opcode=111;
			#100	a=-58173;b=-274485;opcode=111;
			#100	a=-92465;b=560695;opcode=010;
			#100	a=-762901;b=-184522;opcode=100;
			#100	a=-409440;b=-207655;opcode=010;
			#100	a=569368;b=-445231;opcode=111;
			#100	a=-676690;b=-13440;opcode=010;
			#100	a=393129;b=-110342;opcode=110;
			#100	a=612803;b=841863;opcode=111;
			#100	a=65208;b=471091;opcode=001;
			#100	a=380583;b=557785;opcode=001;
			#100	a=264110;b=-272224;opcode=110;
			#100	a=-784102;b=-621832;opcode=000;
			#100	a=-697316;b=-386432;opcode=000;
			#100	a=575651;b=-694871;opcode=110;
			#100	a=779373;b=-998846;opcode=110;
			#100	a=-325857;b=784006;opcode=001;
			#100	a=871599;b=381529;opcode=001;
			#100	a=178695;b=196559;opcode=001;
			#100	a=553557;b=-261096;opcode=000;
			#100	a=-796347;b=-610860;opcode=010;
			#100	a=-247952;b=-160810;opcode=110;
			#100	a=-611927;b=792080;opcode=010;
			#100	a=984386;b=-378809;opcode=001;
			#100	a=-366078;b=-271143;opcode=000;
			#100	a=-980048;b=533775;opcode=000;
			#100	a=-717634;b=182299;opcode=001;
			#100	a=617434;b=765808;opcode=111;
			#100	a=344679;b=-146321;opcode=001;
			#100	a=-885105;b=562735;opcode=000;
			#100	a=258025;b=-84556;opcode=111;
			#100	a=433718;b=64580;opcode=100;
			#100	a=631727;b=648732;opcode=010;
			#100	a=-266474;b=-625896;opcode=000;
			#100	a=-149536;b=879821;opcode=110;
			#100	a=500280;b=-534087;opcode=111;
			#100	a=-193753;b=-354056;opcode=001;
			#100	a=369782;b=-314640;opcode=100;
			#100	a=431668;b=655359;opcode=010;
			#100	a=284639;b=-13436;opcode=001;
			#100	a=-269314;b=-887430;opcode=000;
			#100	a=-206453;b=-207166;opcode=001;
			#100	a=-386068;b=-568021;opcode=111;
			#100	a=330145;b=-985635;opcode=000;
			#100	a=568674;b=-232171;opcode=010;
			#100	a=427259;b=-539841;opcode=110;
			#100	a=426370;b=-245496;opcode=100;
			#100	a=-79420;b=-690843;opcode=001;
			#100	a=905953;b=-789208;opcode=000;
			#100	a=784754;b=29011;opcode=110;
			#100	a=-544283;b=121756;opcode=110;
			#100	a=730655;b=-817730;opcode=100;
			#100	a=287276;b=994018;opcode=010;
			#100	a=-604535;b=-98013;opcode=001;
			#100	a=619792;b=-4848;opcode=001;
			#100	a=56570;b=-870873;opcode=000;
			#100	a=694423;b=-590875;opcode=010;
			#100	a=-294340;b=696458;opcode=110;
			#100	a=348625;b=620885;opcode=001;
			#100	a=-419083;b=-567020;opcode=001;
			#100	a=17344;b=-966129;opcode=001;
			#100	a=-397098;b=839884;opcode=010;
			#100	a=367602;b=-170000;opcode=000;
			#100	a=-246031;b=139853;opcode=000;
			#100	a=-956711;b=-447169;opcode=000;
			#100	a=200417;b=760845;opcode=000;
			#100	a=444782;b=-133056;opcode=000;
			#100	a=300576;b=-500504;opcode=111;
			#100	a=-607883;b=451773;opcode=001;
			#100	a=915324;b=420371;opcode=100;
			#100	a=813999;b=-685799;opcode=010;
			#100	a=-44238;b=907770;opcode=110;
			#100	a=-504388;b=-492975;opcode=000;
			#100	a=715946;b=-114393;opcode=100;
			#100	a=941155;b=-560224;opcode=110;
			#100	a=615820;b=-96234;opcode=001;
			#100	a=461612;b=-901111;opcode=100;
			#100	a=59490;b=62969;opcode=001;
			#100	a=-440687;b=829726;opcode=001;
			#100	a=11623;b=-886390;opcode=010;
			#100	a=-673629;b=253875;opcode=110;
			#100	a=768970;b=945041;opcode=010;
			#100	a=59494;b=139616;opcode=001;
			#100	a=642035;b=-692357;opcode=000;
			#100	a=993861;b=660458;opcode=000;
			#100	a=102233;b=-473374;opcode=110;
			#100	a=-791634;b=49120;opcode=100;
			#100	a=-426906;b=225408;opcode=110;
			#100	a=129786;b=-401977;opcode=001;
			#100	a=858395;b=-950204;opcode=000;
			#100	a=-12611;b=-891249;opcode=100;
			#100	a=-701652;b=699810;opcode=001;
			#100	a=-312983;b=747666;opcode=001;
			#100	a=508388;b=451331;opcode=001;
			#100	a=426801;b=-675408;opcode=110;
			#100	a=313108;b=-867300;opcode=110;
			#100	a=11537;b=-48708;opcode=100;
			#100	a=515988;b=-881999;opcode=110;
			#100	a=-882983;b=462055;opcode=110;
			#100	a=788868;b=448207;opcode=001;
			#100	a=-890868;b=861935;opcode=111;
			#100	a=-27128;b=69675;opcode=110;
			#100	a=-667741;b=-419102;opcode=010;
			#100	a=302619;b=-469703;opcode=001;
			#100	a=-66547;b=424053;opcode=111;
			#100	a=-956273;b=-776381;opcode=010;
			#100	a=-65809;b=-793141;opcode=111;
			#100	a=421230;b=935077;opcode=001;
			#100	a=-227374;b=-744071;opcode=010;
			#100	a=-702718;b=789134;opcode=110;
			#100	a=289272;b=-869179;opcode=100;
			#100	a=417476;b=-214989;opcode=110;
			#100	a=-603001;b=-1155;opcode=110;
			#100	a=-410144;b=-944972;opcode=100;
			#100	a=-556289;b=823663;opcode=000;
			#100	a=-11158;b=404467;opcode=100;
			#100	a=-657343;b=407288;opcode=111;
			#100	a=-129625;b=-15571;opcode=111;
			#100	a=-5548;b=345413;opcode=111;
			#100	a=138385;b=692435;opcode=110;
			#100	a=-813493;b=532912;opcode=100;
			#100	a=416189;b=-486073;opcode=001;
			#100	a=-172108;b=-373708;opcode=010;
			#100	a=404984;b=-17593;opcode=111;
			#100	a=-671023;b=-276328;opcode=000;
			#100	a=31070;b=-166360;opcode=100;
			#100	a=-914398;b=638406;opcode=010;
			#100	a=-672713;b=-434705;opcode=110;
			#100	a=396536;b=774139;opcode=010;
			#100	a=-481791;b=-117675;opcode=111;
			#100	a=50499;b=212196;opcode=010;
			#100	a=578773;b=-894318;opcode=111;
			#100	a=913724;b=873498;opcode=111;
			#100	a=81597;b=-843541;opcode=100;
			#100	a=-636196;b=-178883;opcode=001;
			#100	a=-263742;b=241911;opcode=110;
			#100	a=286564;b=-991505;opcode=001;
			#100	a=-92833;b=-433298;opcode=110;
			#100	a=236786;b=-239610;opcode=111;
			#100	a=993684;b=-948646;opcode=111;
			#100	a=59598;b=-95368;opcode=100;
			#100	a=680542;b=-182507;opcode=001;
			#100	a=-312680;b=-728391;opcode=010;
			#100	a=540975;b=403928;opcode=010;
			#100	a=-383054;b=-189826;opcode=110;
			#100	a=-565591;b=221183;opcode=100;
			#100	a=-967235;b=-849078;opcode=100;
			#100	a=981845;b=-322129;opcode=010;
			#100	a=-987789;b=599319;opcode=000;
			#100	a=-401938;b=-936617;opcode=001;
			#100	a=481294;b=909998;opcode=111;
			#100	a=-827326;b=321060;opcode=001;
			#100	a=421780;b=-515772;opcode=010;
			#100	a=-805971;b=-956353;opcode=100;
			#100	a=-6330;b=-206390;opcode=110;
			#100	a=-532949;b=11751;opcode=111;
			#100	a=-19592;b=-459435;opcode=010;
			#100	a=968386;b=300610;opcode=010;
			#100	a=-536712;b=649172;opcode=001;
			#100	a=-162119;b=-262575;opcode=001;
			#100	a=151633;b=-25947;opcode=111;
			#100	a=536105;b=-816113;opcode=001;
			#100	a=-266094;b=-880766;opcode=010;
			#100	a=393648;b=-188127;opcode=111;
			#100	a=-351982;b=-733685;opcode=000;
			#100	a=-936188;b=-649066;opcode=111;
			#100	a=357612;b=21634;opcode=001;
			#100	a=-29119;b=-356024;opcode=010;
			#100	a=714082;b=177665;opcode=001;
			#100	a=775010;b=242347;opcode=110;
			#100	a=223663;b=111671;opcode=110;
			#100	a=798696;b=916083;opcode=110;
			#100	a=-788593;b=161761;opcode=100;
			#100	a=110757;b=559238;opcode=100;
			#100	a=-420057;b=-761637;opcode=001;
			#100	a=883990;b=645377;opcode=000;
			#100	a=323197;b=109286;opcode=010;
			#100	a=75677;b=-742990;opcode=010;
			#100	a=-670974;b=-562300;opcode=000;
			#100	a=575807;b=141034;opcode=110;
			#100	a=-441437;b=266953;opcode=100;
			#100	a=516962;b=624232;opcode=010;
			#100	a=801228;b=-609270;opcode=001;
			#100	a=-174797;b=527807;opcode=000;
			#100	a=-597089;b=850583;opcode=001;
			#100	a=54878;b=224956;opcode=001;
			#100	a=-349672;b=-201959;opcode=010;
			#100	a=-974298;b=-737326;opcode=111;
			#100	a=-918709;b=-239927;opcode=110;
			#100	a=-246665;b=-150232;opcode=111;
			#100	a=665727;b=-105917;opcode=000;
			#100	a=-263683;b=-207484;opcode=110;
			#100	a=-551365;b=-368506;opcode=000;
			#100	a=127221;b=124911;opcode=111;
			#100	a=661846;b=414440;opcode=001;
			#100	a=716947;b=-779024;opcode=110;
			#100	a=-703461;b=-194179;opcode=001;
			#100	a=-652357;b=48207;opcode=110;
			#100	a=620602;b=524496;opcode=010;
			#100	a=231766;b=837840;opcode=001;
			#100	a=768568;b=188967;opcode=001;
			#100	a=84268;b=-950873;opcode=100;
			#100	a=-111804;b=-852984;opcode=000;
			#100	a=820197;b=342361;opcode=111;
			#100	a=-251684;b=805239;opcode=110;
			#100	a=-895627;b=-964779;opcode=010;
			#100	a=245031;b=817081;opcode=110;
			#100	a=-291219;b=-214430;opcode=010;
			#100	a=373667;b=124676;opcode=000;
			#100	a=-951810;b=-240172;opcode=010;
			#100	a=154687;b=-10090;opcode=010;
			#100	a=284073;b=709783;opcode=001;
			#100	a=549122;b=-727745;opcode=100;
			#100	a=276319;b=411218;opcode=110;
			#100	a=469547;b=26863;opcode=110;
			#100	a=-744110;b=-596775;opcode=010;
			#100	a=194640;b=-246890;opcode=100;
			#100	a=435557;b=583130;opcode=001;
			#100	a=41394;b=760560;opcode=010;
			#100	a=-850712;b=42816;opcode=111;
			#100	a=227365;b=818791;opcode=000;
			#100	a=-535838;b=-585890;opcode=001;
			#100	a=-8280;b=-277637;opcode=000;
			#100	a=-399724;b=-886376;opcode=111;
			#100	a=128738;b=-623686;opcode=110;
			#100	a=-373158;b=-59498;opcode=110;
			#100	a=918705;b=825444;opcode=111;
			#100	a=-509004;b=-674542;opcode=100;
			#100	a=83206;b=806675;opcode=110;
			#100	a=391683;b=816177;opcode=010;
			#100	a=-654367;b=-203184;opcode=110;
			#100	a=-938473;b=210647;opcode=110;
			#100	a=73294;b=-692031;opcode=001;
			#100	a=73619;b=955230;opcode=010;
			#100	a=-750615;b=898668;opcode=000;
			#100	a=-246690;b=174930;opcode=100;
			#100	a=612295;b=417642;opcode=001;
			#100	a=712806;b=615632;opcode=010;
			#100	a=79879;b=-234460;opcode=110;
			#100	a=-499973;b=635614;opcode=010;
			#100	a=776265;b=208392;opcode=000;
			#100	a=781494;b=-408777;opcode=000;
			#100	a=236643;b=-925519;opcode=100;
			#100	a=-89299;b=733155;opcode=100;
			#100	a=-982856;b=-667982;opcode=000;
			#100	a=-367639;b=-308397;opcode=111;
			#100	a=607761;b=-386976;opcode=000;
			#100	a=-956265;b=-178391;opcode=001;
			#100	a=-679503;b=-142552;opcode=110;
			#100	a=609161;b=-280812;opcode=111;
			#100	a=73975;b=96016;opcode=111;
			#100	a=-403056;b=351413;opcode=100;
			#100	a=504654;b=227661;opcode=010;
			#100	a=244619;b=729387;opcode=100;
			#100	a=-921303;b=150489;opcode=100;
			#100	a=844206;b=795211;opcode=010;
			#100	a=657450;b=-793205;opcode=000;
			#100	a=-343908;b=328583;opcode=110;
			#100	a=-255118;b=706328;opcode=111;
			#100	a=475136;b=-669176;opcode=110;
			#100	a=520455;b=910429;opcode=100;
			#100	a=-550033;b=584556;opcode=001;
			#100	a=679435;b=-462358;opcode=110;
			#100	a=-542800;b=-44025;opcode=000;
			#100	a=250584;b=-247314;opcode=111;
			#100	a=-928451;b=-837481;opcode=111;
			#100	a=201247;b=388723;opcode=110;
			#100	a=-653546;b=64206;opcode=010;
			#100	a=-654794;b=-215263;opcode=110;
			#100	a=-430306;b=986995;opcode=100;
			#100	a=341215;b=-575690;opcode=110;
			#100	a=295691;b=338573;opcode=000;
			#100	a=-166309;b=-981369;opcode=000;
			#100	a=34918;b=-841318;opcode=000;
			#100	a=-818734;b=32927;opcode=110;
			#100	a=-596759;b=-757130;opcode=100;
			#100	a=-476819;b=871002;opcode=000;
			#100	a=-566888;b=-455509;opcode=010;
			#100	a=-48010;b=-876858;opcode=010;
			#100	a=-685144;b=782267;opcode=100;
			#100	a=-134533;b=-555780;opcode=100;
			#100	a=895072;b=455591;opcode=001;
			#100	a=-310392;b=-758412;opcode=111;
			#100	a=458421;b=466364;opcode=100;
			#100	a=18768;b=-640213;opcode=010;
			#100	a=732123;b=802440;opcode=111;
			#100	a=-875614;b=-857384;opcode=100;
			#100	a=274483;b=217416;opcode=001;
			#100	a=-476273;b=623207;opcode=001;
			#100	a=59113;b=-4242;opcode=001;
			#100	a=415626;b=-84730;opcode=110;
			#100	a=891735;b=352306;opcode=100;
			#100	a=-863899;b=-377941;opcode=100;
			#100	a=216928;b=209078;opcode=100;
			#100	a=-120527;b=-218586;opcode=110;
			#100	a=542665;b=7176;opcode=001;
			#100	a=275198;b=-407840;opcode=110;
			#100	a=521701;b=712812;opcode=111;
			#100	a=-519827;b=-56966;opcode=100;
			#100	a=909930;b=-256715;opcode=110;
			#100	a=-119907;b=723279;opcode=111;
			#100	a=550913;b=-885889;opcode=111;
			#100	a=520566;b=886439;opcode=111;
			#100	a=447293;b=-880609;opcode=010;
			#100	a=-113437;b=-300646;opcode=100;
			#100	a=-281287;b=984876;opcode=010;
			#100	a=991082;b=-930012;opcode=010;
			#100	a=499376;b=263885;opcode=000;
			#100	a=-579433;b=-317894;opcode=100;
			#100	a=-918660;b=-689773;opcode=010;
			#100	a=-502059;b=986655;opcode=001;
			#100	a=-480367;b=-485831;opcode=010;
			#100	a=524843;b=33453;opcode=110;
			#100	a=985370;b=-906056;opcode=111;
			#100	a=754870;b=525263;opcode=000;
			#100	a=732307;b=-671907;opcode=100;
			#100	a=531648;b=-596962;opcode=010;
			#100	a=-298970;b=-687648;opcode=100;
			#100	a=-622531;b=136453;opcode=001;
			#100	a=217193;b=-490845;opcode=111;
			#100	a=-549712;b=376637;opcode=000;
			#100	a=305452;b=-345419;opcode=000;
			#100	a=807579;b=-780812;opcode=111;
			#100	a=83735;b=-350988;opcode=001;
			#100	a=-683903;b=494073;opcode=111;
			#100	a=-45983;b=603260;opcode=111;
			#100	a=488805;b=86434;opcode=100;
			#100	a=393592;b=179146;opcode=110;
			#100	a=-82452;b=895634;opcode=010;
			#100	a=-661469;b=235688;opcode=111;
			#100	a=15645;b=-637160;opcode=111;
			#100	a=-506662;b=699577;opcode=100;
			#100	a=-456886;b=-184639;opcode=110;
			#100	a=810629;b=-448656;opcode=010;
			#100	a=-138466;b=-683647;opcode=001;
			#100	a=308835;b=246931;opcode=000;
			#100	a=812340;b=675684;opcode=110;
			#100	a=995159;b=-249683;opcode=111;
			#100	a=590188;b=884103;opcode=000;
			#100	a=-88621;b=-952010;opcode=001;
			#100	a=694191;b=943140;opcode=000;
			#100	a=839718;b=-213519;opcode=000;
			#100	a=-216964;b=299859;opcode=010;
			#100	a=-878351;b=799689;opcode=100;
			#100	a=6660;b=989517;opcode=010;
			#100	a=-441382;b=958167;opcode=100;
			#100	a=584095;b=-69777;opcode=010;
			#100	a=-487246;b=61737;opcode=110;
			#100	a=-769187;b=307674;opcode=111;
			#100	a=676337;b=-365987;opcode=000;
			#100	a=-852492;b=-104230;opcode=010;
			#100	a=-410116;b=657110;opcode=010;
			#100	a=-282194;b=896576;opcode=100;
			#100	a=445470;b=-740359;opcode=111;
			#100	a=-479935;b=330530;opcode=111;
			#100	a=631212;b=928826;opcode=110;
			#100	a=-300962;b=241174;opcode=110;
			#100	a=-361267;b=263002;opcode=000;
			#100	a=-497740;b=-780837;opcode=111;
			#100	a=295841;b=16229;opcode=110;
			#100	a=621800;b=22817;opcode=000;
			#100	a=-372392;b=820279;opcode=110;
			#100	a=894506;b=503804;opcode=000;
			#100	a=-390865;b=-135243;opcode=000;
			#100	a=644359;b=33182;opcode=110;
			#100	a=-123388;b=535183;opcode=111;
			#100	a=-660255;b=861607;opcode=100;
			#100	a=13739;b=236286;opcode=001;
			#100	a=965223;b=-356819;opcode=111;
			#100	a=418753;b=-87985;opcode=001;
			#100	a=-20663;b=733625;opcode=111;
			#100	a=-160046;b=99005;opcode=111;
			#100	a=150794;b=74663;opcode=110;
			#100	a=-736564;b=703854;opcode=001;
			#100	a=734149;b=-759305;opcode=111;
			#100	a=913900;b=-786233;opcode=001;
			#100	a=-120066;b=-601914;opcode=111;
			#100	a=-776774;b=608377;opcode=000;
			#100	a=448457;b=649696;opcode=100;
			#100	a=-127339;b=-472874;opcode=110;
			#100	a=209318;b=169995;opcode=000;
			#100	a=929008;b=902464;opcode=001;
			#100	a=-809583;b=273758;opcode=110;
			#100	a=-281411;b=9197;opcode=001;
			#100	a=-872641;b=-58101;opcode=000;
			#100	a=226336;b=688026;opcode=010;
			#100	a=861291;b=-811707;opcode=001;
			#100	a=-454551;b=218322;opcode=100;
			#100	a=-454181;b=32345;opcode=100;
			#100	a=563698;b=-496756;opcode=010;
			#100	a=936592;b=519341;opcode=100;
			#100	a=-682712;b=-684388;opcode=001;
			#100	a=367074;b=-535444;opcode=010;
			#100	a=497530;b=-764519;opcode=110;
			#100	a=926789;b=862229;opcode=100;
			#100	a=918836;b=-822108;opcode=111;
			#100	a=492703;b=656614;opcode=001;
			#100	a=-855695;b=-718319;opcode=111;
			#100	a=622043;b=-729611;opcode=111;
			#100	a=-453802;b=-637666;opcode=111;
			#100	a=-171904;b=138141;opcode=110;
			#100	a=-443853;b=501200;opcode=110;
			#100	a=300301;b=289507;opcode=110;
			#100	a=-11047;b=607863;opcode=001;
			#100	a=-182340;b=685936;opcode=100;
			#100	a=763394;b=-255786;opcode=000;
			#100	a=-23692;b=-580905;opcode=100;
			#100	a=769733;b=-985588;opcode=000;
			#100	a=-579781;b=-82624;opcode=001;
			#100	a=-281777;b=377309;opcode=000;
			#100	a=625006;b=44014;opcode=001;
			#100	a=304631;b=-508105;opcode=111;
			#100	a=-382998;b=495643;opcode=100;
			#100	a=133974;b=-589958;opcode=000;
			#100	a=212266;b=-823940;opcode=010;
			#100	a=59129;b=-709850;opcode=110;
			#100	a=-477253;b=-682967;opcode=000;
			#100	a=168779;b=316286;opcode=001;
			#100	a=-546679;b=191701;opcode=000;
			#100	a=387334;b=304755;opcode=100;
			#100	a=1153;b=-662423;opcode=100;
			#100	a=527689;b=427621;opcode=000;
			#100	a=655804;b=807776;opcode=010;
			#100	a=662749;b=343006;opcode=110;
			#100	a=-487743;b=400907;opcode=010;
			#100	a=-441031;b=-324174;opcode=110;
			#100	a=-245483;b=57391;opcode=100;
			#100	a=-52414;b=-766983;opcode=110;
			#100	a=-623391;b=-373345;opcode=110;
			#100	a=-550254;b=-187237;opcode=100;

		end
endmodule

